library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_0 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"31",X"F0",X"4F",X"E7",X"C3",X"B4",X"01",X"FF",X"AF",X"77",X"23",X"10",X"FC",X"C9",X"FF",X"FF",
		X"D5",X"07",X"5F",X"16",X"00",X"19",X"D1",X"C9",X"E1",X"18",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AF",X"32",X"00",X"50",X"32",X"C0",X"50",X"C9",X"E7",X"3E",X"01",X"32",X"00",X"50",X"C9",X"FF",
		X"18",X"1C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CD",X"AA",X"01",X"0F",X"0F",X"0F",X"E6",X"1E",
		X"5F",X"16",X"00",X"21",X"CB",X"01",X"19",X"5E",X"23",X"56",X"EB",X"F1",X"F5",X"E9",X"CB",X"27",
		X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"EB",X"E9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"ED",X"73",X"1E",X"48",X"31",X"C0",X"4F",X"08",X"D9",X"E7",
		X"DD",X"E5",X"FD",X"E5",X"CD",X"DD",X"01",X"FD",X"E1",X"DD",X"E1",X"0E",X"03",X"21",X"B0",X"4B",
		X"06",X"08",X"11",X"06",X"00",X"7E",X"FE",X"01",X"23",X"20",X"1B",X"79",X"A6",X"23",X"28",X"03",
		X"35",X"28",X"0C",X"19",X"10",X"EF",X"EF",X"D9",X"08",X"ED",X"7B",X"1E",X"48",X"ED",X"45",X"2B",
		X"CB",X"FE",X"2B",X"36",X"03",X"23",X"23",X"18",X"EA",X"31",X"F0",X"4F",X"FB",X"0E",X"00",X"21",
		X"B0",X"4B",X"06",X"08",X"11",X"08",X"00",X"7E",X"CB",X"7F",X"20",X"04",X"FE",X"02",X"30",X"06",
		X"0C",X"19",X"10",X"F3",X"18",X"E7",X"F3",X"79",X"32",X"00",X"48",X"7E",X"36",X"02",X"23",X"CB",
		X"BE",X"23",X"36",X"00",X"23",X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"23",X"EB",X"FE",X"04",
		X"20",X"04",X"50",X"59",X"FB",X"E9",X"F9",X"FE",X"02",X"28",X"04",X"1A",X"C1",X"18",X"01",X"F1",
		X"C1",X"D1",X"E1",X"FD",X"E1",X"DD",X"E1",X"FB",X"C9",X"CD",X"9A",X"01",X"36",X"04",X"23",X"72",
		X"23",X"72",X"23",X"71",X"23",X"70",X"18",X"E7",X"CD",X"9A",X"01",X"72",X"18",X"E1",X"CD",X"97",
		X"01",X"7E",X"FE",X"02",X"C2",X"A9",X"00",X"23",X"7E",X"CB",X"7F",X"20",X"15",X"E6",X"40",X"4F",
		X"F1",X"F5",X"E6",X"0F",X"B1",X"77",X"23",X"70",X"2B",X"2B",X"36",X"01",X"CD",X"89",X"01",X"C3",
		X"A9",X"00",X"CB",X"BE",X"1E",X"06",X"19",X"7E",X"18",X"B2",X"CD",X"9A",X"01",X"CB",X"BE",X"7E",
		X"B7",X"28",X"AC",X"FE",X"04",X"28",X"A8",X"1E",X"07",X"19",X"70",X"11",X"FA",X"FF",X"19",X"CB",
		X"F6",X"CB",X"FE",X"FE",X"01",X"20",X"98",X"2B",X"36",X"03",X"18",X"93",X"CD",X"9A",X"01",X"7E",
		X"B7",X"28",X"8C",X"CB",X"FE",X"18",X"88",X"CD",X"97",X"01",X"72",X"C3",X"A9",X"00",X"CD",X"9A",
		X"01",X"1E",X"05",X"19",X"71",X"23",X"70",X"C3",X"EF",X"00",X"CD",X"97",X"01",X"23",X"CB",X"76",
		X"CB",X"B6",X"1E",X"06",X"19",X"7E",X"C3",X"EC",X"00",X"01",X"03",X"00",X"09",X"EB",X"21",X"02",
		X"00",X"39",X"EB",X"73",X"23",X"72",X"C9",X"3A",X"00",X"48",X"E6",X"0F",X"21",X"B0",X"4B",X"16",
		X"00",X"5F",X"CB",X"23",X"CB",X"23",X"CB",X"23",X"19",X"C9",X"DD",X"E3",X"FD",X"E5",X"E5",X"D5",
		X"C5",X"F5",X"DD",X"E9",X"21",X"00",X"48",X"01",X"00",X"18",X"36",X"00",X"23",X"0B",X"78",X"B1",
		X"20",X"F8",X"3E",X"07",X"01",X"30",X"35",X"FF",X"C3",X"A9",X"00",X"F9",X"00",X"08",X"01",X"0E",
		X"01",X"0E",X"01",X"3A",X"01",X"5C",X"01",X"67",X"01",X"6E",X"01",X"7A",X"01",X"3A",X"C0",X"50",
		X"2F",X"32",X"20",X"48",X"21",X"80",X"50",X"36",X"01",X"36",X"00",X"21",X"03",X"48",X"3A",X"00",
		X"50",X"2F",X"E6",X"A0",X"20",X"07",X"7E",X"B7",X"20",X"12",X"C3",X"80",X"02",X"36",X"06",X"FE",
		X"80",X"CA",X"80",X"02",X"3E",X"01",X"32",X"07",X"50",X"C3",X"80",X"02",X"AF",X"32",X"07",X"50",
		X"36",X"00",X"23",X"7E",X"3C",X"77",X"23",X"86",X"B7",X"28",X"36",X"CB",X"7F",X"20",X"32",X"47",
		X"AF",X"32",X"04",X"48",X"23",X"7E",X"80",X"77",X"FE",X"64",X"30",X"1A",X"05",X"CB",X"20",X"48",
		X"06",X"00",X"21",X"41",X"02",X"09",X"11",X"08",X"48",X"06",X"02",X"CD",X"54",X"3D",X"18",X"11",
		X"00",X"01",X"00",X"02",X"00",X"03",X"3E",X"63",X"32",X"06",X"48",X"21",X"09",X"09",X"22",X"07",
		X"48",X"21",X"02",X"48",X"CB",X"7E",X"20",X"1B",X"E5",X"21",X"49",X"42",X"DD",X"21",X"07",X"48",
		X"1E",X"0B",X"06",X"02",X"0E",X"00",X"CD",X"8A",X"3D",X"3E",X"08",X"16",X"00",X"1E",X"00",X"CD",
		X"20",X"2C",X"E1",X"2B",X"CB",X"7E",X"CB",X"FE",X"20",X"06",X"3E",X"07",X"01",X"35",X"35",X"FF",
		X"21",X"88",X"4B",X"DD",X"21",X"F0",X"4F",X"FD",X"21",X"60",X"50",X"06",X"08",X"CB",X"7E",X"20",
		X"4F",X"4E",X"0C",X"3A",X"21",X"48",X"57",X"CB",X"FE",X"23",X"7E",X"CB",X"42",X"28",X"09",X"EE",
		X"C0",X"E6",X"C0",X"5F",X"3E",X"3F",X"A6",X"B3",X"07",X"07",X"DD",X"77",X"00",X"23",X"7E",X"CB",
		X"42",X"28",X"04",X"ED",X"44",X"C6",X"10",X"D6",X"02",X"FD",X"77",X"00",X"23",X"7E",X"DD",X"77",
		X"01",X"23",X"7E",X"CB",X"42",X"28",X"04",X"ED",X"44",X"C6",X"10",X"FD",X"77",X"01",X"23",X"DD",
		X"23",X"DD",X"23",X"FD",X"23",X"FD",X"23",X"05",X"CA",X"5E",X"2D",X"0D",X"28",X"AF",X"18",X"B3",
		X"11",X"05",X"00",X"19",X"DD",X"23",X"DD",X"23",X"FD",X"23",X"FD",X"23",X"10",X"9F",X"C3",X"5E",
		X"2D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E5",X"D1",X"06",X"D2",X"CF",X"21",X"4B",X"03",X"3A",X"02",X"48",X"CB",X"77",X"20",X"0C",X"CD",
		X"4D",X"0E",X"D5",X"21",X"33",X"03",X"CD",X"E1",X"3D",X"EB",X"D1",X"4E",X"23",X"06",X"01",X"7E",
		X"FE",X"FF",X"C8",X"FE",X"C0",X"38",X"05",X"E6",X"3F",X"47",X"23",X"7E",X"12",X"13",X"10",X"FC",
		X"23",X"18",X"EA",X"C1",X"03",X"62",X"04",X"2E",X"05",X"00",X"06",X"CF",X"06",X"A1",X"07",X"71",
		X"08",X"45",X"09",X"13",X"0A",X"E7",X"0A",X"B6",X"0B",X"88",X"0C",X"64",X"D0",X"00",X"11",X"25",
		X"35",X"45",X"15",X"25",X"35",X"43",X"C3",X"00",X"10",X"C3",X"00",X"46",X"C6",X"00",X"16",X"C3",
		X"00",X"21",X"C3",X"00",X"36",X"C6",X"00",X"26",X"C3",X"00",X"32",X"C3",X"00",X"26",X"C6",X"00",
		X"36",X"C3",X"00",X"43",X"C3",X"00",X"16",X"C6",X"00",X"46",X"00",X"27",X"00",X"14",X"C3",X"00",
		X"46",X"C6",X"00",X"16",X"C3",X"00",X"25",X"C3",X"00",X"36",X"C6",X"00",X"26",X"00",X"47",X"00",
		X"36",X"C3",X"00",X"26",X"C6",X"00",X"36",X"C3",X"00",X"47",X"C3",X"00",X"16",X"C6",X"00",X"46",
		X"C3",X"00",X"18",X"C3",X"00",X"46",X"C6",X"00",X"16",X"C3",X"00",X"29",X"C3",X"00",X"36",X"C6",
		X"00",X"26",X"00",X"57",X"00",X"3A",X"C3",X"00",X"22",X"15",X"45",X"35",X"25",X"15",X"45",X"34",
		X"FF",X"1E",X"C4",X"00",X"01",X"47",X"05",X"55",X"05",X"17",X"03",X"C8",X"00",X"06",X"02",X"07",
		X"05",X"07",X"04",X"06",X"C8",X"00",X"3A",X"05",X"0B",X"05",X"0B",X"35",X"09",X"C8",X"00",X"06",
		X"01",X"08",X"25",X"08",X"03",X"26",X"C4",X"00",X"01",X"07",X"25",X"05",X"0B",X"0B",X"07",X"05",
		X"15",X"0B",X"0B",X"07",X"15",X"05",X"03",X"06",X"06",X"01",X"07",X"09",X"26",X"0A",X"07",X"03",
		X"06",X"46",X"06",X"01",X"07",X"09",X"06",X"36",X"C6",X"06",X"26",X"0A",X"09",X"C3",X"06",X"46",
		X"16",X"06",X"06",X"46",X"0A",X"09",X"C4",X"06",X"16",X"06",X"36",X"06",X"06",X"0A",X"08",X"04",
		X"26",X"06",X"06",X"02",X"08",X"09",X"06",X"0A",X"08",X"24",X"06",X"06",X"42",X"05",X"15",X"08",
		X"0B",X"3B",X"05",X"05",X"48",X"0B",X"0B",X"05",X"05",X"08",X"04",X"C4",X"00",X"06",X"02",X"07",
		X"05",X"07",X"04",X"06",X"C8",X"00",X"1A",X"05",X"0B",X"15",X"0B",X"05",X"39",X"C8",X"00",X"06",
		X"01",X"08",X"05",X"08",X"03",X"06",X"C8",X"00",X"02",X"08",X"05",X"55",X"05",X"48",X"04",X"C8",
		X"00",X"FF",X"33",X"01",X"05",X"35",X"05",X"03",X"21",X"05",X"05",X"55",X"03",X"21",X"05",X"05",
		X"35",X"43",X"0A",X"07",X"17",X"05",X"0B",X"08",X"47",X"15",X"07",X"08",X"08",X"05",X"07",X"07",
		X"09",X"06",X"06",X"0A",X"07",X"09",X"01",X"0B",X"05",X"0B",X"33",X"70",X"01",X"09",X"46",X"06",
		X"26",X"C4",X"06",X"46",X"02",X"05",X"04",X"1A",X"47",X"09",X"36",X"16",X"06",X"02",X"0B",X"0B",
		X"18",X"09",X"06",X"01",X"35",X"03",X"06",X"0A",X"08",X"0B",X"0B",X"04",X"01",X"39",X"0A",X"25",
		X"08",X"0B",X"0B",X"07",X"0B",X"0B",X"08",X"35",X"09",X"1A",X"03",X"06",X"06",X"0A",X"05",X"35",
		X"09",X"06",X"06",X"46",X"2A",X"05",X"05",X"09",X"26",X"06",X"06",X"46",X"0A",X"05",X"05",X"09",
		X"C3",X"06",X"0A",X"05",X"45",X"09",X"06",X"06",X"02",X"09",X"3A",X"25",X"07",X"0B",X"0B",X"08",
		X"0B",X"0B",X"07",X"05",X"09",X"0A",X"04",X"01",X"1B",X"0B",X"07",X"09",X"16",X"22",X"05",X"04",
		X"16",X"3A",X"07",X"0B",X"0B",X"13",X"C3",X"06",X"0A",X"08",X"39",X"01",X"05",X"13",X"C6",X"06",
		X"56",X"06",X"0A",X"44",X"70",X"02",X"0B",X"05",X"0B",X"04",X"0A",X"08",X"39",X"36",X"26",X"0A",
		X"08",X"08",X"05",X"07",X"07",X"08",X"45",X"28",X"57",X"0B",X"15",X"08",X"08",X"09",X"02",X"05",
		X"05",X"15",X"04",X"02",X"15",X"05",X"05",X"04",X"02",X"05",X"25",X"05",X"04",X"FF",X"35",X"01",
		X"05",X"15",X"27",X"05",X"05",X"07",X"05",X"57",X"05",X"45",X"07",X"B5",X"35",X"23",X"0A",X"07",
		X"05",X"0B",X"05",X"45",X"0B",X"35",X"0B",X"25",X"05",X"0B",X"05",X"47",X"09",X"06",X"36",X"70",
		X"1A",X"07",X"05",X"09",X"70",X"0A",X"05",X"37",X"09",X"70",X"06",X"06",X"0A",X"0B",X"07",X"0B",
		X"0B",X"25",X"0B",X"05",X"0B",X"05",X"0B",X"0B",X"07",X"0B",X"09",X"56",X"06",X"36",X"06",X"06",
		X"41",X"0B",X"15",X"0B",X"03",X"46",X"06",X"16",X"06",X"46",X"26",X"06",X"06",X"0A",X"04",X"36",
		X"0A",X"05",X"09",X"06",X"02",X"09",X"C3",X"06",X"02",X"08",X"0B",X"08",X"25",X"0B",X"0B",X"05",
		X"3B",X"0B",X"15",X"08",X"0B",X"08",X"24",X"01",X"07",X"4B",X"07",X"05",X"0B",X"0B",X"05",X"0B",
		X"0B",X"45",X"07",X"0B",X"07",X"43",X"06",X"06",X"16",X"0A",X"03",X"06",X"3A",X"05",X"19",X"06",
		X"01",X"09",X"36",X"06",X"06",X"16",X"36",X"C3",X"06",X"02",X"0B",X"05",X"0B",X"24",X"06",X"16",
		X"06",X"06",X"06",X"2A",X"0B",X"08",X"0B",X"3B",X"45",X"0B",X"05",X"0B",X"05",X"0B",X"0B",X"28",
		X"0B",X"09",X"06",X"46",X"70",X"0A",X"08",X"05",X"09",X"70",X"0A",X"15",X"38",X"09",X"70",X"06",
		X"06",X"0A",X"08",X"05",X"0B",X"15",X"05",X"0B",X"35",X"0B",X"25",X"05",X"0B",X"45",X"08",X"29",
		X"02",X"05",X"05",X"48",X"05",X"15",X"08",X"05",X"58",X"05",X"05",X"08",X"05",X"05",X"04",X"FF",
		X"37",X"01",X"05",X"27",X"05",X"07",X"07",X"35",X"03",X"70",X"01",X"07",X"05",X"55",X"05",X"13",
		X"0A",X"05",X"08",X"33",X"06",X"02",X"05",X"08",X"03",X"06",X"0A",X"27",X"05",X"33",X"06",X"0A",
		X"45",X"03",X"0A",X"0B",X"45",X"17",X"35",X"08",X"04",X"46",X"0A",X"05",X"08",X"09",X"0A",X"05",
		X"3B",X"04",X"0A",X"07",X"0B",X"07",X"35",X"05",X"09",X"0A",X"05",X"15",X"09",X"0A",X"05",X"0B",
		X"05",X"09",X"16",X"36",X"16",X"01",X"05",X"0B",X"0B",X"25",X"03",X"06",X"1A",X"A5",X"08",X"25",
		X"09",X"36",X"06",X"02",X"0B",X"45",X"09",X"06",X"70",X"0A",X"09",X"2A",X"05",X"05",X"07",X"08",
		X"49",X"0A",X"05",X"0B",X"35",X"29",X"02",X"17",X"04",X"46",X"0A",X"05",X"45",X"09",X"70",X"0A",
		X"08",X"47",X"0B",X"05",X"4B",X"05",X"0B",X"05",X"09",X"5A",X"07",X"13",X"0A",X"07",X"0B",X"03",
		X"06",X"02",X"05",X"0B",X"07",X"0B",X"35",X"04",X"C3",X"06",X"16",X"06",X"36",X"26",X"0A",X"05",
		X"15",X"09",X"36",X"36",X"01",X"03",X"4A",X"C6",X"0B",X"08",X"57",X"07",X"09",X"06",X"16",X"06",
		X"06",X"06",X"12",X"0B",X"09",X"06",X"16",X"06",X"70",X"06",X"36",X"0A",X"08",X"0B",X"0B",X"19",
		X"0A",X"05",X"04",X"26",X"46",X"02",X"0B",X"05",X"09",X"06",X"0A",X"25",X"0B",X"04",X"06",X"02",
		X"05",X"05",X"08",X"08",X"05",X"38",X"B5",X"48",X"08",X"18",X"05",X"38",X"05",X"04",X"FF",X"3C",
		X"01",X"05",X"07",X"17",X"05",X"05",X"37",X"07",X"05",X"15",X"07",X"07",X"35",X"95",X"13",X"0A",
		X"05",X"3B",X"0B",X"05",X"45",X"09",X"06",X"01",X"25",X"09",X"36",X"01",X"27",X"09",X"0A",X"05",
		X"09",X"2A",X"07",X"05",X"2B",X"08",X"5B",X"07",X"0B",X"08",X"2B",X"0B",X"09",X"0A",X"05",X"14",
		X"06",X"0A",X"07",X"0B",X"03",X"06",X"16",X"06",X"70",X"06",X"16",X"36",X"0A",X"05",X"27",X"08",
		X"34",X"06",X"36",X"0A",X"4B",X"04",X"0A",X"07",X"0B",X"08",X"09",X"0A",X"05",X"08",X"03",X"41",
		X"08",X"09",X"06",X"02",X"25",X"09",X"06",X"02",X"35",X"09",X"1A",X"05",X"55",X"0B",X"0B",X"05",
		X"0B",X"08",X"17",X"05",X"4B",X"08",X"05",X"07",X"19",X"0A",X"25",X"05",X"04",X"0A",X"35",X"09",
		X"70",X"0A",X"05",X"3B",X"05",X"47",X"09",X"06",X"0A",X"15",X"07",X"45",X"0B",X"25",X"08",X"07",
		X"2B",X"07",X"0B",X"05",X"09",X"06",X"06",X"0A",X"05",X"0B",X"35",X"0B",X"B5",X"33",X"06",X"16",
		X"06",X"06",X"01",X"08",X"0B",X"09",X"2A",X"05",X"29",X"70",X"0A",X"05",X"C4",X"0B",X"4B",X"0B",
		X"03",X"36",X"06",X"06",X"41",X"0B",X"05",X"0B",X"07",X"39",X"26",X"06",X"26",X"56",X"1A",X"08",
		X"08",X"19",X"06",X"06",X"0A",X"05",X"39",X"06",X"0A",X"0B",X"18",X"08",X"09",X"02",X"25",X"03",
		X"06",X"02",X"08",X"08",X"15",X"08",X"08",X"28",X"08",X"25",X"05",X"48",X"05",X"A5",X"18",X"04",
		X"FF",X"3F",X"01",X"17",X"05",X"27",X"05",X"35",X"07",X"07",X"57",X"05",X"15",X"07",X"05",X"37",
		X"13",X"06",X"06",X"01",X"1B",X"35",X"45",X"09",X"26",X"0A",X"05",X"45",X"0B",X"03",X"06",X"06",
		X"0A",X"08",X"0B",X"0B",X"05",X"07",X"08",X"0B",X"38",X"07",X"B5",X"0B",X"0B",X"48",X"09",X"0A",
		X"07",X"0B",X"3B",X"15",X"09",X"70",X"06",X"70",X"0A",X"35",X"4B",X"0B",X"37",X"09",X"0A",X"39",
		X"02",X"2B",X"07",X"08",X"27",X"08",X"07",X"08",X"07",X"0B",X"04",X"0A",X"09",X"0A",X"0B",X"07",
		X"09",X"3A",X"07",X"0B",X"07",X"0B",X"23",X"06",X"4A",X"07",X"3B",X"49",X"96",X"56",X"36",X"C4",
		X"06",X"16",X"06",X"06",X"4A",X"19",X"26",X"06",X"06",X"36",X"06",X"06",X"2A",X"19",X"C3",X"06",
		X"26",X"16",X"C3",X"06",X"16",X"06",X"0A",X"2B",X"08",X"19",X"06",X"42",X"0B",X"28",X"0B",X"48",
		X"09",X"1A",X"08",X"0B",X"09",X"0A",X"09",X"01",X"0B",X"28",X"07",X"08",X"07",X"08",X"27",X"08",
		X"1B",X"03",X"2A",X"09",X"0A",X"38",X"0B",X"4B",X"05",X"09",X"70",X"06",X"70",X"0A",X"05",X"0B",
		X"0B",X"08",X"09",X"0A",X"07",X"0B",X"0B",X"05",X"08",X"17",X"0B",X"07",X"08",X"05",X"2B",X"0B",
		X"07",X"49",X"16",X"06",X"02",X"2B",X"35",X"05",X"09",X"06",X"0A",X"A5",X"15",X"0B",X"04",X"06",
		X"06",X"02",X"08",X"05",X"28",X"05",X"05",X"58",X"08",X"18",X"05",X"45",X"08",X"05",X"18",X"04",
		X"FF",X"47",X"01",X"07",X"07",X"07",X"37",X"05",X"07",X"15",X"07",X"47",X"A5",X"27",X"05",X"07",
		X"43",X"06",X"26",X"06",X"46",X"0A",X"05",X"4B",X"05",X"3B",X"0B",X"07",X"0B",X"05",X"39",X"06",
		X"3A",X"18",X"0B",X"08",X"0B",X"35",X"0B",X"05",X"09",X"56",X"06",X"16",X"21",X"08",X"09",X"0A",
		X"25",X"09",X"70",X"0A",X"05",X"0B",X"15",X"0B",X"48",X"0B",X"0B",X"0B",X"05",X"19",X"4A",X"05",
		X"08",X"07",X"18",X"07",X"2B",X"05",X"0B",X"05",X"0B",X"48",X"0B",X"05",X"39",X"0A",X"47",X"15",
		X"0B",X"05",X"4B",X"0B",X"45",X"09",X"70",X"0A",X"07",X"48",X"07",X"09",X"0A",X"0B",X"05",X"0B",
		X"13",X"06",X"0A",X"07",X"08",X"27",X"08",X"1B",X"05",X"3B",X"09",X"1A",X"08",X"55",X"0B",X"0B",
		X"38",X"09",X"1A",X"05",X"4B",X"35",X"0B",X"33",X"06",X"06",X"0A",X"27",X"05",X"4B",X"09",X"70",
		X"0A",X"2B",X"05",X"3B",X"B5",X"2B",X"0B",X"0B",X"09",X"96",X"3A",X"05",X"0B",X"0B",X"07",X"04",
		X"0A",X"05",X"0B",X"07",X"08",X"0B",X"44",X"06",X"3A",X"0B",X"03",X"26",X"46",X"0A",X"05",X"0B",
		X"15",X"0B",X"49",X"70",X"0A",X"35",X"09",X"06",X"22",X"0B",X"0B",X"08",X"0B",X"07",X"4B",X"07",
		X"09",X"0A",X"37",X"0B",X"07",X"49",X"2A",X"05",X"09",X"1A",X"35",X"09",X"36",X"06",X"06",X"3A",
		X"09",X"56",X"16",X"06",X"06",X"02",X"05",X"08",X"38",X"05",X"18",X"08",X"28",X"18",X"08",X"28",
		X"08",X"08",X"38",X"04",X"FF",X"3F",X"01",X"15",X"05",X"07",X"55",X"47",X"07",X"07",X"A5",X"07",
		X"47",X"35",X"07",X"45",X"13",X"06",X"01",X"05",X"0B",X"05",X"09",X"06",X"16",X"01",X"08",X"0B",
		X"07",X"09",X"21",X"09",X"0A",X"0B",X"35",X"0B",X"05",X"0B",X"18",X"28",X"0B",X"33",X"16",X"26",
		X"0A",X"09",X"06",X"16",X"0A",X"05",X"09",X"70",X"0A",X"05",X"05",X"09",X"06",X"46",X"16",X"36",
		X"06",X"56",X"2A",X"3B",X"17",X"0B",X"37",X"08",X"37",X"17",X"C4",X"0B",X"08",X"08",X"09",X"C3",
		X"06",X"0A",X"0B",X"25",X"0B",X"0B",X"09",X"06",X"36",X"0A",X"05",X"07",X"09",X"02",X"C3",X"0B",
		X"08",X"07",X"09",X"06",X"1A",X"49",X"16",X"0A",X"45",X"0B",X"14",X"70",X"36",X"26",X"06",X"01",
		X"29",X"0A",X"09",X"36",X"0A",X"08",X"09",X"70",X"0A",X"43",X"01",X"1B",X"C4",X"0B",X"18",X"08",
		X"0B",X"0B",X"25",X"0B",X"07",X"08",X"09",X"96",X"36",X"06",X"36",X"42",X"0B",X"15",X"45",X"2B",
		X"08",X"B5",X"09",X"4A",X"05",X"09",X"0A",X"08",X"0B",X"0B",X"07",X"38",X"07",X"07",X"0B",X"07",
		X"47",X"0B",X"0B",X"07",X"09",X"2A",X"05",X"09",X"06",X"06",X"70",X"06",X"06",X"16",X"06",X"16",
		X"26",X"06",X"06",X"16",X"0A",X"05",X"0B",X"29",X"0A",X"37",X"08",X"0B",X"4B",X"0B",X"0B",X"3B",
		X"18",X"09",X"06",X"02",X"05",X"08",X"58",X"08",X"08",X"05",X"08",X"38",X"34",X"02",X"08",X"05",
		X"08",X"04",X"FF",X"4A",X"01",X"07",X"07",X"07",X"B5",X"45",X"37",X"05",X"07",X"45",X"07",X"15",
		X"07",X"05",X"13",X"0A",X"0B",X"19",X"0A",X"05",X"07",X"2B",X"07",X"18",X"07",X"08",X"07",X"5B",
		X"23",X"06",X"36",X"22",X"3B",X"08",X"27",X"0B",X"0B",X"29",X"70",X"0A",X"47",X"0B",X"0B",X"1B",
		X"29",X"0A",X"05",X"4B",X"03",X"56",X"06",X"16",X"0A",X"07",X"09",X"0A",X"09",X"36",X"06",X"06",
		X"0A",X"03",X"06",X"0A",X"0B",X"09",X"36",X"2A",X"0B",X"49",X"06",X"3A",X"1B",X"09",X"06",X"1A",
		X"0B",X"49",X"36",X"06",X"0A",X"0B",X"04",X"0A",X"28",X"1B",X"09",X"06",X"3A",X"49",X"06",X"0A",
		X"08",X"0B",X"4B",X"08",X"0B",X"05",X"0B",X"35",X"09",X"0A",X"08",X"09",X"06",X"0A",X"09",X"70",
		X"2A",X"1B",X"37",X"0B",X"47",X"0B",X"25",X"0B",X"09",X"70",X"0A",X"39",X"36",X"0A",X"07",X"09",
		X"A6",X"0A",X"0B",X"3B",X"09",X"01",X"09",X"0A",X"27",X"09",X"06",X"16",X"46",X"36",X"0A",X"08",
		X"09",X"46",X"06",X"3A",X"29",X"0A",X"08",X"09",X"4A",X"09",X"02",X"0B",X"0B",X"0B",X"25",X"0B",
		X"0B",X"0B",X"08",X"0B",X"0B",X"25",X"0B",X"08",X"09",X"01",X"09",X"32",X"0B",X"07",X"5B",X"0B",
		X"19",X"70",X"0A",X"0B",X"35",X"0B",X"03",X"36",X"0A",X"28",X"07",X"04",X"2A",X"04",X"36",X"22",
		X"07",X"44",X"3A",X"07",X"08",X"1B",X"49",X"02",X"05",X"48",X"05",X"28",X"45",X"08",X"95",X"18",
		X"05",X"28",X"48",X"35",X"08",X"04",X"FF",X"4E",X"01",X"05",X"27",X"95",X"17",X"07",X"35",X"07",
		X"27",X"05",X"17",X"05",X"07",X"35",X"43",X"06",X"70",X"0A",X"35",X"2B",X"4B",X"23",X"1A",X"0B",
		X"35",X"0B",X"55",X"09",X"70",X"06",X"0A",X"07",X"08",X"07",X"09",X"0A",X"0B",X"09",X"0A",X"23",
		X"06",X"01",X"08",X"17",X"29",X"3A",X"5B",X"03",X"06",X"06",X"16",X"06",X"46",X"16",X"0A",X"4B",
		X"09",X"31",X"0B",X"19",X"06",X"02",X"1B",X"3B",X"0B",X"0B",X"3B",X"0B",X"3B",X"2B",X"C3",X"0B",
		X"04",X"06",X"1A",X"07",X"0B",X"09",X"42",X"0B",X"0B",X"08",X"0B",X"0B",X"04",X"2A",X"0B",X"37",
		X"09",X"96",X"36",X"26",X"3A",X"05",X"2B",X"09",X"70",X"0A",X"1B",X"05",X"09",X"16",X"06",X"26",
		X"06",X"0A",X"0B",X"0B",X"07",X"0B",X"0B",X"17",X"0B",X"0B",X"43",X"1A",X"0B",X"39",X"06",X"4A",
		X"08",X"29",X"06",X"36",X"06",X"46",X"A6",X"06",X"26",X"0A",X"09",X"4A",X"28",X"09",X"36",X"01",
		X"4B",X"0B",X"2B",X"C4",X"0B",X"4B",X"C3",X"0B",X"03",X"06",X"1A",X"3B",X"04",X"C3",X"06",X"0A",
		X"39",X"0A",X"0B",X"09",X"B6",X"42",X"0B",X"09",X"0A",X"08",X"07",X"08",X"29",X"0A",X"4B",X"08",
		X"0B",X"14",X"3A",X"28",X"07",X"38",X"19",X"06",X"70",X"2A",X"35",X"0B",X"58",X"09",X"01",X"2B",
		X"05",X"1B",X"05",X"09",X"70",X"06",X"02",X"05",X"18",X"05",X"28",X"05",X"18",X"04",X"42",X"05",
		X"08",X"25",X"08",X"05",X"24",X"FF",X"49",X"01",X"05",X"07",X"27",X"37",X"95",X"07",X"05",X"37",
		X"05",X"07",X"45",X"07",X"35",X"03",X"0A",X"17",X"0B",X"4B",X"08",X"07",X"29",X"70",X"0A",X"47",
		X"08",X"37",X"09",X"11",X"29",X"0A",X"4B",X"09",X"36",X"11",X"38",X"0B",X"07",X"0B",X"08",X"07",
		X"09",X"2A",X"0B",X"09",X"36",X"0A",X"08",X"0B",X"09",X"01",X"0B",X"14",X"5A",X"07",X"19",X"0A",
		X"08",X"09",X"46",X"0A",X"09",X"70",X"2A",X"0B",X"0B",X"3B",X"07",X"0B",X"2B",X"0B",X"09",X"70",
		X"0A",X"09",X"1A",X"08",X"07",X"09",X"06",X"26",X"06",X"46",X"36",X"06",X"36",X"0A",X"17",X"38",
		X"09",X"26",X"70",X"4A",X"0B",X"1B",X"C3",X"0B",X"2B",X"C3",X"0B",X"09",X"70",X"06",X"3A",X"07",
		X"08",X"09",X"26",X"46",X"06",X"16",X"06",X"A6",X"46",X"0A",X"28",X"17",X"09",X"0A",X"09",X"70",
		X"0A",X"0B",X"0B",X"0B",X"38",X"1B",X"4B",X"0B",X"09",X"70",X"0A",X"09",X"B6",X"3A",X"07",X"0B",
		X"59",X"12",X"0B",X"03",X"3A",X"08",X"09",X"0A",X"17",X"09",X"06",X"4A",X"0B",X"19",X"06",X"0A",
		X"25",X"39",X"0A",X"29",X"01",X"2B",X"09",X"36",X"4A",X"09",X"06",X"16",X"4A",X"0B",X"3B",X"B5",
		X"4B",X"08",X"0B",X"1B",X"04",X"0A",X"0B",X"0B",X"09",X"0A",X"08",X"0B",X"08",X"2B",X"15",X"09",
		X"70",X"0A",X"08",X"07",X"58",X"09",X"02",X"19",X"02",X"05",X"28",X"05",X"18",X"05",X"08",X"25",
		X"08",X"35",X"08",X"05",X"08",X"25",X"04",X"FF",X"43",X"01",X"05",X"07",X"05",X"47",X"07",X"15",
		X"07",X"35",X"03",X"01",X"35",X"07",X"45",X"03",X"4A",X"B5",X"0B",X"33",X"0A",X"09",X"01",X"5B",
		X"03",X"4A",X"09",X"01",X"0B",X"05",X"19",X"36",X"01",X"08",X"0B",X"24",X"4A",X"39",X"06",X"1A",
		X"29",X"02",X"1B",X"08",X"33",X"96",X"0A",X"19",X"01",X"08",X"07",X"08",X"09",X"46",X"0A",X"08",
		X"47",X"08",X"03",X"0A",X"09",X"0A",X"08",X"0B",X"17",X"09",X"70",X"4A",X"2B",X"09",X"70",X"0A",
		X"27",X"0B",X"58",X"09",X"0A",X"03",X"26",X"0A",X"08",X"07",X"0B",X"08",X"0B",X"07",X"04",X"46",
		X"36",X"01",X"09",X"0A",X"3B",X"0B",X"4B",X"05",X"3B",X"09",X"70",X"0A",X"2B",X"35",X"0B",X"0B",
		X"0B",X"19",X"4A",X"04",X"06",X"0A",X"07",X"08",X"3B",X"07",X"0B",X"08",X"03",X"26",X"06",X"22",
		X"09",X"0A",X"05",X"1B",X"38",X"09",X"70",X"0A",X"1B",X"09",X"70",X"0A",X"08",X"0B",X"15",X"09",
		X"16",X"01",X"08",X"07",X"08",X"07",X"39",X"96",X"2A",X"07",X"0B",X"07",X"38",X"03",X"06",X"0A",
		X"09",X"31",X"0B",X"57",X"09",X"46",X"36",X"06",X"06",X"0A",X"0B",X"23",X"4A",X"09",X"3A",X"0B",
		X"0B",X"04",X"16",X"06",X"0A",X"0B",X"38",X"0B",X"39",X"02",X"0B",X"0B",X"09",X"06",X"06",X"42",
		X"07",X"08",X"0B",X"09",X"0A",X"05",X"09",X"22",X"07",X"04",X"36",X"06",X"02",X"08",X"05",X"28",
		X"05",X"38",X"08",X"48",X"05",X"28",X"05",X"18",X"A5",X"18",X"24",X"FF",X"DD",X"21",X"41",X"40",
		X"FD",X"21",X"30",X"48",X"01",X"0E",X"0F",X"C5",X"DD",X"E5",X"C5",X"FD",X"7E",X"00",X"B7",X"28",
		X"3B",X"47",X"E6",X"F0",X"FE",X"70",X"28",X"1D",X"FE",X"90",X"38",X"28",X"CD",X"4B",X"0F",X"78",
		X"E6",X"0F",X"FE",X"06",X"3E",X"1C",X"28",X"02",X"3E",X"18",X"DD",X"E5",X"E1",X"01",X"02",X"02",
		X"CD",X"1E",X"3D",X"18",X"17",X"DD",X"E5",X"E1",X"3E",X"C0",X"1E",X"17",X"01",X"02",X"02",X"CD",
		X"1E",X"3D",X"18",X"08",X"78",X"DD",X"E5",X"CD",X"41",X"0E",X"DD",X"E1",X"C1",X"DD",X"23",X"DD",
		X"23",X"FD",X"23",X"10",X"B5",X"3E",X"23",X"06",X"02",X"FF",X"DD",X"E1",X"01",X"40",X"00",X"DD",
		X"09",X"C1",X"0D",X"20",X"A2",X"CD",X"4D",X"0E",X"FE",X"00",X"C0",X"DD",X"21",X"FB",X"0F",X"21",
		X"62",X"40",X"CD",X"1D",X"0E",X"DD",X"21",X"FB",X"0F",X"21",X"78",X"40",X"CD",X"1D",X"0E",X"DD",
		X"21",X"04",X"10",X"21",X"E2",X"42",X"CD",X"1D",X"0E",X"DD",X"21",X"04",X"10",X"21",X"F8",X"42",
		X"CD",X"1D",X"0E",X"21",X"A4",X"40",X"1E",X"02",X"CD",X"14",X"0E",X"21",X"BA",X"40",X"1E",X"01",
		X"CD",X"14",X"0E",X"21",X"24",X"43",X"1E",X"03",X"CD",X"14",X"0E",X"21",X"3A",X"43",X"1E",X"04",
		X"CD",X"14",X"0E",X"C9",X"3E",X"C4",X"01",X"02",X"02",X"CD",X"1E",X"3D",X"C9",X"01",X"03",X"03",
		X"1E",X"17",X"C5",X"E5",X"C5",X"E5",X"DD",X"7E",X"00",X"01",X"02",X"02",X"CD",X"1E",X"3D",X"DD",
		X"23",X"E1",X"23",X"23",X"C1",X"10",X"ED",X"E1",X"01",X"40",X"00",X"09",X"C1",X"0D",X"20",X"E2",
		X"C9",X"DD",X"E5",X"E1",X"1E",X"03",X"DD",X"21",X"77",X"89",X"C3",X"39",X"0F",X"3A",X"E7",X"49",
		X"FE",X"0C",X"D8",X"D6",X"0C",X"18",X"F9",X"21",X"D4",X"0E",X"22",X"14",X"4A",X"21",X"41",X"40",
		X"FD",X"21",X"30",X"48",X"01",X"0E",X"0F",X"C5",X"E5",X"C5",X"E5",X"FD",X"7E",X"00",X"47",X"E6",
		X"F0",X"28",X"1D",X"FE",X"70",X"30",X"19",X"E5",X"2A",X"14",X"4A",X"7E",X"21",X"CC",X"0E",X"CD",
		X"E1",X"3D",X"D5",X"DD",X"E1",X"78",X"E6",X"F0",X"CD",X"4B",X"0F",X"E1",X"78",X"CD",X"50",X"89",
		X"E1",X"23",X"23",X"FD",X"23",X"C1",X"10",X"D1",X"E1",X"01",X"40",X"00",X"09",X"C1",X"0D",X"20",
		X"C6",X"2A",X"14",X"4A",X"5E",X"21",X"E5",X"0E",X"16",X"00",X"19",X"7E",X"16",X"00",X"1E",X"00",
		X"CD",X"20",X"2C",X"3E",X"23",X"06",X"08",X"FF",X"2A",X"14",X"4A",X"23",X"22",X"14",X"4A",X"7E",
		X"FE",X"FF",X"20",X"99",X"3E",X"01",X"CD",X"8E",X"2C",X"C3",X"E9",X"0E",X"77",X"89",X"A3",X"89",
		X"CF",X"89",X"27",X"8A",X"00",X"01",X"02",X"01",X"00",X"01",X"02",X"01",X"00",X"01",X"02",X"02",
		X"01",X"02",X"01",X"02",X"FF",X"01",X"02",X"03",X"02",X"DD",X"21",X"41",X"40",X"FD",X"21",X"30",
		X"48",X"01",X"0E",X"0F",X"C5",X"DD",X"E5",X"C5",X"FD",X"7E",X"00",X"B7",X"DD",X"E5",X"C4",X"18",
		X"0F",X"DD",X"E1",X"C1",X"DD",X"23",X"DD",X"23",X"FD",X"23",X"10",X"EB",X"DD",X"E1",X"01",X"40",
		X"00",X"DD",X"09",X"C1",X"0D",X"20",X"DD",X"C9",X"47",X"E6",X"F0",X"C8",X"FE",X"80",X"20",X"07",
		X"78",X"E6",X"0F",X"FD",X"77",X"00",X"C9",X"FE",X"50",X"28",X"12",X"FE",X"50",X"D0",X"CD",X"4B",
		X"0F",X"78",X"DD",X"E5",X"E1",X"DD",X"21",X"27",X"8A",X"CD",X"50",X"89",X"C9",X"DD",X"E5",X"E1",
		X"3E",X"D0",X"1E",X"05",X"01",X"02",X"02",X"CD",X"1E",X"3D",X"C9",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"3D",X"21",X"5D",X"0F",X"16",X"00",X"5F",X"19",X"5E",X"C9",X"01",X"02",X"03",
		X"04",X"07",X"06",X"17",X"00",X"5B",X"5C",X"5D",X"7D",X"4D",X"E6",X"C0",X"6F",X"B7",X"11",X"40",
		X"40",X"ED",X"52",X"38",X"26",X"29",X"29",X"7C",X"FE",X"0E",X"30",X"1F",X"6F",X"87",X"87",X"87",
		X"87",X"95",X"6F",X"79",X"E6",X"1F",X"FE",X"1E",X"30",X"11",X"CB",X"47",X"28",X"0D",X"3D",X"CB",
		X"3F",X"85",X"5F",X"16",X"00",X"21",X"30",X"48",X"19",X"7E",X"C9",X"3E",X"FF",X"C9",X"7C",X"E6",
		X"F0",X"D6",X"20",X"38",X"F6",X"FE",X"D1",X"30",X"F2",X"67",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"4F",X"7C",X"91",X"67",X"7D",X"ED",X"44",X"E6",X"F8",X"D6",X"08",X"38",X"DC",X"FE",
		X"E1",X"30",X"D8",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"84",X"C3",X"92",X"0F",X"11",
		X"30",X"48",X"B7",X"ED",X"52",X"7D",X"26",X"20",X"FE",X"0F",X"38",X"0A",X"D6",X"0F",X"47",X"7C",
		X"C6",X"10",X"67",X"78",X"18",X"F2",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"C6",X"08",
		X"ED",X"44",X"6F",X"C9",X"CD",X"CF",X"0F",X"CD",X"BC",X"3D",X"C9",X"C0",X"C0",X"C0",X"C0",X"00",
		X"C0",X"C0",X"00",X"C0",X"C0",X"00",X"C0",X"C0",X"00",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"FF",
		X"31",X"60",X"4F",X"21",X"14",X"4A",X"06",X"38",X"CF",X"21",X"BE",X"24",X"22",X"40",X"4A",X"AF",
		X"32",X"42",X"4A",X"FD",X"21",X"14",X"4A",X"3A",X"E6",X"49",X"47",X"05",X"CD",X"EF",X"3E",X"21",
		X"22",X"27",X"11",X"14",X"4A",X"01",X"24",X"00",X"ED",X"B0",X"CD",X"97",X"1A",X"06",X"03",X"C5",
		X"CD",X"90",X"11",X"3E",X"23",X"06",X"18",X"FF",X"21",X"88",X"4B",X"06",X"19",X"CF",X"3E",X"23",
		X"06",X"0C",X"FF",X"C1",X"10",X"E9",X"3E",X"23",X"06",X"01",X"FF",X"3E",X"45",X"FF",X"3E",X"02",
		X"01",X"50",X"8C",X"FF",X"3E",X"01",X"01",X"78",X"86",X"FF",X"3E",X"03",X"01",X"48",X"3F",X"FF",
		X"3A",X"DA",X"49",X"CB",X"47",X"16",X"00",X"28",X"02",X"16",X"FF",X"1E",X"00",X"3E",X"00",X"CD",
		X"20",X"2C",X"3E",X"23",X"06",X"01",X"FF",X"21",X"E4",X"49",X"35",X"20",X"55",X"EB",X"21",X"28",
		X"25",X"3A",X"E7",X"49",X"FE",X"0A",X"38",X"02",X"3E",X"0A",X"06",X"00",X"4F",X"09",X"7E",X"EB",
		X"77",X"21",X"E1",X"49",X"35",X"F5",X"3A",X"DA",X"49",X"CB",X"47",X"20",X"21",X"7E",X"FE",X"18",
		X"20",X"1C",X"3A",X"DA",X"49",X"CB",X"47",X"CB",X"C7",X"32",X"DA",X"49",X"3E",X"09",X"16",X"00",
		X"1E",X"00",X"CD",X"20",X"2C",X"3E",X"00",X"16",X"FF",X"1E",X"00",X"CD",X"20",X"2C",X"CD",X"12",
		X"3F",X"F1",X"20",X"0E",X"3A",X"02",X"48",X"CB",X"4F",X"CB",X"CF",X"32",X"02",X"48",X"FD",X"36",
		X"11",X"20",X"FD",X"21",X"14",X"4A",X"3A",X"01",X"48",X"CB",X"67",X"28",X"2A",X"FD",X"6E",X"24",
		X"FD",X"66",X"25",X"2B",X"FD",X"75",X"24",X"FD",X"74",X"25",X"7C",X"B5",X"20",X"19",X"FD",X"6E",
		X"26",X"FD",X"66",X"27",X"FD",X"7E",X"29",X"77",X"3A",X"01",X"48",X"CB",X"67",X"CB",X"A7",X"32",
		X"01",X"48",X"3E",X"0D",X"CD",X"8E",X"2C",X"FD",X"7E",X"08",X"FE",X"04",X"28",X"0E",X"FE",X"03",
		X"28",X"0A",X"3A",X"01",X"48",X"CB",X"4F",X"20",X"03",X"CD",X"61",X"1B",X"FD",X"7E",X"09",X"21",
		X"35",X"11",X"F7",X"18",X"0A",X"DE",X"11",X"DE",X"11",X"02",X"16",X"1D",X"16",X"57",X"16",X"FD",
		X"7E",X"08",X"21",X"F7",X"11",X"F7",X"FD",X"7E",X"30",X"B7",X"28",X"3E",X"FE",X"01",X"20",X"2D",
		X"FD",X"7E",X"32",X"B7",X"28",X"05",X"FD",X"35",X"32",X"18",X"2F",X"FD",X"7E",X"1B",X"FE",X"36",
		X"20",X"12",X"FD",X"36",X"30",X"02",X"FD",X"36",X"31",X"40",X"FD",X"36",X"1B",X"25",X"FD",X"36",
		X"1D",X"4F",X"18",X"16",X"FD",X"34",X"1B",X"FD",X"36",X"32",X"08",X"18",X"0D",X"FD",X"35",X"31",
		X"20",X"08",X"FD",X"36",X"1B",X"00",X"FD",X"36",X"30",X"00",X"CD",X"90",X"11",X"C3",X"82",X"10",
		X"21",X"18",X"4A",X"11",X"8E",X"4B",X"01",X"04",X"00",X"ED",X"B0",X"21",X"34",X"4A",X"11",X"93",
		X"4B",X"01",X"04",X"00",X"ED",X"B0",X"21",X"2F",X"4A",X"11",X"9D",X"4B",X"01",X"04",X"00",X"ED",
		X"B0",X"FD",X"7E",X"09",X"FE",X"03",X"28",X"27",X"21",X"2B",X"4A",X"11",X"98",X"4B",X"01",X"04",
		X"00",X"ED",X"B0",X"21",X"14",X"4A",X"11",X"89",X"4B",X"01",X"04",X"00",X"ED",X"B0",X"AF",X"32",
		X"88",X"4B",X"32",X"8D",X"4B",X"32",X"92",X"4B",X"32",X"97",X"4B",X"32",X"9C",X"4B",X"C9",X"21",
		X"14",X"4A",X"11",X"98",X"4B",X"01",X"04",X"00",X"ED",X"B0",X"21",X"2B",X"4A",X"11",X"89",X"4B",
		X"01",X"04",X"00",X"ED",X"B0",X"18",X"D7",X"03",X"12",X"68",X"14",X"E7",X"17",X"8C",X"14",X"32",
		X"18",X"B2",X"15",X"CD",X"B2",X"1A",X"FD",X"7E",X"08",X"FE",X"05",X"28",X"33",X"CD",X"BC",X"19",
		X"20",X"2E",X"FD",X"66",X"21",X"FD",X"6E",X"23",X"CD",X"9E",X"0F",X"E6",X"F0",X"FE",X"80",X"20",
		X"1F",X"FD",X"7E",X"08",X"FE",X"01",X"28",X"18",X"3E",X"11",X"CD",X"8E",X"2C",X"3E",X"05",X"16",
		X"00",X"1E",X"00",X"CD",X"20",X"2C",X"FD",X"36",X"08",X"05",X"FD",X"7E",X"0E",X"FD",X"77",X"11",
		X"3A",X"01",X"48",X"CB",X"4F",X"28",X"20",X"CD",X"BC",X"19",X"C2",X"05",X"14",X"3E",X"00",X"CD",
		X"8E",X"2C",X"3A",X"01",X"48",X"CB",X"5F",X"C2",X"A6",X"19",X"3E",X"23",X"06",X"40",X"FF",X"3E",
		X"47",X"06",X"10",X"FF",X"C3",X"A6",X"19",X"3A",X"02",X"48",X"CB",X"4F",X"28",X"1C",X"FD",X"7E",
		X"11",X"B7",X"CA",X"9C",X"19",X"FD",X"35",X"11",X"CD",X"BC",X"19",X"20",X"0A",X"CD",X"F2",X"19",
		X"E6",X"F0",X"28",X"03",X"C3",X"9C",X"19",X"AF",X"18",X"03",X"CD",X"FE",X"1A",X"CB",X"67",X"CA",
		X"20",X"13",X"47",X"FD",X"7E",X"08",X"FE",X"05",X"78",X"CA",X"24",X"13",X"47",X"3E",X"03",X"FD",
		X"BE",X"09",X"78",X"CA",X"24",X"13",X"FD",X"CB",X"1F",X"46",X"C2",X"24",X"13",X"FD",X"CB",X"01",
		X"46",X"C2",X"24",X"13",X"FD",X"CB",X"03",X"46",X"C2",X"24",X"13",X"3A",X"E2",X"49",X"3C",X"32",
		X"E2",X"49",X"FD",X"36",X"0A",X"03",X"CD",X"87",X"1A",X"FD",X"36",X"1F",X"01",X"FD",X"36",X"08",
		X"03",X"FD",X"CB",X"0E",X"46",X"20",X"16",X"FD",X"7E",X"03",X"E6",X"0F",X"0E",X"20",X"FD",X"CB",
		X"0E",X"4E",X"20",X"03",X"81",X"18",X"17",X"ED",X"44",X"E6",X"0F",X"18",X"F7",X"FD",X"7E",X"01",
		X"C6",X"08",X"E6",X"0F",X"0E",X"20",X"FD",X"CB",X"0E",X"4E",X"28",X"EB",X"18",X"E6",X"FD",X"77",
		X"12",X"FD",X"36",X"13",X"00",X"21",X"8D",X"26",X"CD",X"1B",X"1A",X"21",X"16",X"27",X"CD",X"5E",
		X"1A",X"3E",X"04",X"CD",X"8E",X"2C",X"3E",X"07",X"16",X"00",X"1E",X"00",X"CD",X"20",X"2C",X"C9",
		X"FD",X"36",X"1F",X"00",X"CD",X"CA",X"19",X"FD",X"77",X"0F",X"5F",X"FE",X"04",X"20",X"1D",X"FD",
		X"7E",X"2F",X"B7",X"28",X"05",X"FD",X"35",X"2F",X"18",X"16",X"FD",X"7E",X"0A",X"FE",X"02",X"28",
		X"4B",X"FD",X"36",X"0A",X"02",X"D5",X"CD",X"87",X"1A",X"D1",X"18",X"40",X"FD",X"36",X"2F",X"0C",
		X"7B",X"EE",X"02",X"FD",X"BE",X"0E",X"20",X"1D",X"FD",X"7E",X"08",X"FE",X"05",X"20",X"05",X"FD",
		X"5E",X"0E",X"18",X"11",X"FD",X"36",X"0A",X"06",X"D5",X"CD",X"87",X"1A",X"D1",X"CD",X"BC",X"19",
		X"C2",X"D3",X"13",X"18",X"26",X"7B",X"FD",X"BE",X"0E",X"20",X"11",X"FD",X"36",X"0A",X"06",X"D5",
		X"CD",X"87",X"1A",X"D1",X"CD",X"BC",X"19",X"C2",X"05",X"14",X"18",X"0F",X"CD",X"BC",X"19",X"C2",
		X"05",X"14",X"7B",X"FE",X"04",X"20",X"04",X"FD",X"7E",X"0E",X"5F",X"D5",X"CD",X"89",X"17",X"D1",
		X"7B",X"CD",X"EB",X"3D",X"A6",X"C2",X"D3",X"13",X"FD",X"7E",X"0E",X"5F",X"CD",X"EB",X"3D",X"A6",
		X"C2",X"D3",X"13",X"7B",X"D6",X"01",X"E6",X"03",X"5F",X"CD",X"EB",X"3D",X"A6",X"20",X"04",X"7B",
		X"EE",X"02",X"5F",X"FD",X"7E",X"0A",X"FE",X"02",X"28",X"09",X"FD",X"36",X"0A",X"02",X"D5",X"CD",
		X"87",X"1A",X"D1",X"FD",X"73",X"0F",X"FD",X"7E",X"0F",X"FD",X"BE",X"0E",X"CA",X"05",X"14",X"3E",
		X"05",X"CD",X"8E",X"2C",X"FD",X"36",X"08",X"01",X"FD",X"36",X"10",X"04",X"FD",X"4E",X"0F",X"FD",
		X"7E",X"0E",X"FD",X"71",X"0E",X"21",X"A2",X"26",X"CD",X"E1",X"3D",X"EB",X"CD",X"5E",X"1A",X"21",
		X"DA",X"26",X"CD",X"1B",X"1A",X"FD",X"7E",X"08",X"FE",X"05",X"28",X"04",X"CD",X"06",X"1A",X"D0",
		X"21",X"32",X"25",X"FD",X"7E",X"08",X"FE",X"05",X"20",X"03",X"21",X"3A",X"25",X"FD",X"7E",X"0E",
		X"CD",X"E1",X"3D",X"D5",X"C1",X"FD",X"66",X"01",X"FD",X"6E",X"03",X"CD",X"83",X"3D",X"FD",X"74",
		X"01",X"FD",X"75",X"03",X"FD",X"66",X"05",X"FD",X"6E",X"07",X"CD",X"83",X"3D",X"FD",X"74",X"05",
		X"FD",X"75",X"07",X"FD",X"66",X"21",X"FD",X"6E",X"23",X"CD",X"83",X"3D",X"FD",X"74",X"21",X"FD",
		X"75",X"23",X"FD",X"7E",X"09",X"FE",X"03",X"C0",X"FD",X"66",X"18",X"FD",X"6E",X"1A",X"CD",X"83",
		X"3D",X"FD",X"74",X"18",X"FD",X"75",X"1A",X"C9",X"FD",X"7E",X"10",X"B7",X"28",X"06",X"FD",X"35",
		X"10",X"C3",X"06",X"12",X"CD",X"7A",X"14",X"C3",X"06",X"12",X"FD",X"36",X"08",X"00",X"21",X"FA",
		X"26",X"CD",X"5E",X"1A",X"CD",X"97",X"1A",X"FD",X"CB",X"10",X"BE",X"C9",X"CD",X"06",X"1A",X"D0",
		X"FD",X"7E",X"12",X"B7",X"CA",X"0D",X"15",X"21",X"0A",X"27",X"FD",X"7E",X"13",X"FE",X"08",X"28",
		X"0A",X"FD",X"7E",X"12",X"21",X"16",X"27",X"FE",X"08",X"20",X"03",X"CD",X"5E",X"1A",X"FD",X"7E",
		X"13",X"0E",X"02",X"FE",X"08",X"38",X"0F",X"0E",X"01",X"FE",X"18",X"38",X"09",X"FD",X"7E",X"12",
		X"FE",X"09",X"30",X"02",X"0E",X"02",X"FD",X"7E",X"12",X"91",X"30",X"01",X"AF",X"FD",X"77",X"12",
		X"79",X"FD",X"86",X"13",X"FD",X"77",X"13",X"C5",X"CD",X"98",X"17",X"C1",X"79",X"FD",X"CB",X"0E",
		X"46",X"20",X"15",X"FD",X"CB",X"0E",X"4E",X"20",X"01",X"ED",X"44",X"FD",X"86",X"03",X"FD",X"77",
		X"03",X"FD",X"77",X"07",X"FD",X"77",X"23",X"C9",X"FD",X"CB",X"0E",X"4E",X"28",X"01",X"ED",X"44",
		X"FD",X"86",X"01",X"FD",X"77",X"01",X"FD",X"77",X"05",X"FD",X"77",X"21",X"C9",X"3E",X"07",X"CD",
		X"8E",X"2C",X"FD",X"36",X"08",X"00",X"FD",X"36",X"09",X"00",X"FD",X"36",X"28",X"00",X"FD",X"36",
		X"0A",X"06",X"CD",X"87",X"1A",X"21",X"14",X"4A",X"11",X"2B",X"4A",X"01",X"08",X"00",X"ED",X"B0",
		X"AF",X"32",X"2B",X"4A",X"32",X"2F",X"4A",X"21",X"DA",X"26",X"CD",X"1B",X"1A",X"21",X"FA",X"26",
		X"CD",X"5E",X"1A",X"FD",X"7E",X"0E",X"CD",X"E0",X"19",X"CD",X"9E",X"0F",X"FE",X"FF",X"28",X"5C",
		X"E6",X"F0",X"28",X"58",X"FE",X"80",X"CA",X"21",X"12",X"FE",X"90",X"D2",X"AC",X"1C",X"FE",X"70",
		X"20",X"03",X"C3",X"6C",X"17",X"FD",X"36",X"08",X"02",X"47",X"C5",X"CD",X"D5",X"17",X"C1",X"28",
		X"2A",X"78",X"21",X"42",X"25",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"3D",X"16",X"00",
		X"5F",X"19",X"7E",X"FD",X"77",X"19",X"FD",X"77",X"1D",X"FD",X"36",X"09",X"01",X"FD",X"36",X"16",
		X"00",X"3E",X"0C",X"16",X"00",X"1E",X"00",X"CD",X"20",X"2C",X"C9",X"FD",X"66",X"21",X"FD",X"6E",
		X"23",X"CD",X"9E",X"0F",X"E5",X"CD",X"F4",X"0F",X"D1",X"CD",X"CD",X"1B",X"CD",X"FE",X"1A",X"C3",
		X"24",X"13",X"FD",X"7E",X"10",X"CB",X"BF",X"B7",X"28",X"06",X"FD",X"35",X"10",X"C3",X"06",X"12",
		X"3E",X"02",X"FD",X"B6",X"10",X"FD",X"77",X"10",X"FD",X"CB",X"10",X"7E",X"FD",X"CB",X"10",X"BE",
		X"20",X"2B",X"FD",X"CB",X"10",X"FE",X"FD",X"4E",X"11",X"79",X"C6",X"01",X"FE",X"04",X"38",X"01",
		X"AF",X"FD",X"77",X"11",X"C5",X"21",X"DA",X"26",X"CD",X"1E",X"1A",X"C1",X"79",X"21",X"A2",X"26",
		X"CD",X"E1",X"3D",X"EB",X"FD",X"7E",X"11",X"CD",X"61",X"1A",X"C3",X"06",X"12",X"21",X"FA",X"26",
		X"18",X"F2",X"FD",X"36",X"09",X"03",X"21",X"FA",X"26",X"CD",X"5E",X"1A",X"CD",X"97",X"1A",X"FD",
		X"CB",X"10",X"BE",X"21",X"DA",X"26",X"CD",X"1B",X"1A",X"FD",X"36",X"19",X"1A",X"3A",X"01",X"48",
		X"CB",X"7F",X"C8",X"CD",X"FE",X"1A",X"CB",X"67",X"C8",X"FD",X"36",X"1F",X"01",X"FD",X"36",X"09",
		X"04",X"FD",X"7E",X"08",X"FE",X"05",X"FD",X"7E",X"0E",X"20",X"03",X"FD",X"7E",X"11",X"FD",X"77",
		X"2A",X"FD",X"36",X"2B",X"02",X"21",X"18",X"25",X"CD",X"E1",X"3D",X"FD",X"73",X"17",X"3E",X"0F",
		X"16",X"00",X"1E",X"00",X"CD",X"20",X"2C",X"FD",X"7E",X"2B",X"FD",X"35",X"2B",X"20",X"1D",X"FD",
		X"36",X"2B",X"02",X"FD",X"7E",X"2A",X"21",X"18",X"25",X"CD",X"E1",X"3D",X"FD",X"7E",X"17",X"B7",
		X"28",X"07",X"7B",X"FD",X"BE",X"17",X"20",X"01",X"7A",X"FD",X"77",X"17",X"FD",X"66",X"18",X"FD",
		X"6E",X"1A",X"FD",X"CB",X"2A",X"46",X"28",X"0D",X"7C",X"FE",X"F8",X"D2",X"5D",X"17",X"FE",X"08",
		X"DA",X"5D",X"17",X"18",X"1B",X"7D",X"FD",X"CB",X"2A",X"4E",X"20",X"07",X"FE",X"10",X"DA",X"5D",
		X"17",X"18",X"0D",X"FE",X"20",X"30",X"09",X"FE",X"18",X"D2",X"5D",X"17",X"FD",X"36",X"17",X"00",
		X"FD",X"CB",X"2A",X"46",X"20",X"1F",X"7D",X"C6",X"08",X"6F",X"E6",X"0F",X"FE",X"01",X"38",X"45",
		X"FE",X"0E",X"30",X"41",X"7D",X"E6",X"F0",X"0E",X"E8",X"FD",X"CB",X"2A",X"4E",X"20",X"02",X"0E",
		X"08",X"81",X"6F",X"18",X"0F",X"7C",X"E6",X"0F",X"FE",X"01",X"38",X"29",X"FE",X"0E",X"30",X"25",
		X"7C",X"E6",X"F0",X"67",X"E5",X"CD",X"9E",X"0F",X"D1",X"FE",X"FF",X"28",X"18",X"E6",X"F0",X"28",
		X"14",X"FE",X"80",X"28",X"10",X"FE",X"70",X"28",X"0C",X"FE",X"90",X"30",X"23",X"E5",X"CD",X"F4",
		X"0F",X"D1",X"CD",X"CD",X"1B",X"21",X"20",X"25",X"FD",X"7E",X"2A",X"CD",X"E1",X"3D",X"D5",X"C1",
		X"FD",X"66",X"18",X"FD",X"6E",X"1A",X"CD",X"83",X"3D",X"FD",X"74",X"18",X"FD",X"75",X"1A",X"C9",
		X"FD",X"36",X"30",X"01",X"FD",X"36",X"32",X"08",X"FD",X"36",X"1B",X"34",X"FD",X"36",X"1D",X"49",
		X"FD",X"72",X"1C",X"FD",X"73",X"1E",X"CD",X"4A",X"17",X"21",X"6B",X"17",X"CD",X"04",X"3E",X"3E",
		X"11",X"16",X"00",X"1E",X"00",X"CD",X"20",X"2C",X"18",X"BB",X"7E",X"E6",X"0F",X"77",X"F5",X"CD",
		X"F4",X"0F",X"F1",X"DD",X"21",X"77",X"89",X"1E",X"01",X"CD",X"50",X"89",X"C9",X"FD",X"36",X"17",
		X"00",X"FD",X"36",X"09",X"00",X"C9",X"00",X"00",X"01",X"00",X"00",X"00",X"3A",X"01",X"48",X"CB",
		X"57",X"CB",X"D7",X"32",X"01",X"48",X"FD",X"36",X"08",X"04",X"3E",X"00",X"CD",X"8E",X"2C",X"3E",
		X"0B",X"16",X"00",X"1E",X"00",X"CD",X"20",X"2C",X"C9",X"FD",X"66",X"21",X"FD",X"6E",X"23",X"CD",
		X"9E",X"0F",X"E6",X"0F",X"CD",X"D8",X"19",X"C9",X"CD",X"D5",X"17",X"C0",X"CD",X"89",X"17",X"FD",
		X"7E",X"0E",X"D6",X"01",X"E6",X"03",X"5F",X"CD",X"EB",X"3D",X"A6",X"20",X"04",X"7B",X"EE",X"02",
		X"5F",X"FD",X"73",X"0E",X"21",X"16",X"27",X"FD",X"7E",X"13",X"FE",X"08",X"38",X"0D",X"21",X"0A",
		X"27",X"FD",X"7E",X"12",X"FE",X"09",X"30",X"03",X"21",X"16",X"27",X"CD",X"5E",X"1A",X"21",X"8D",
		X"26",X"CD",X"1B",X"1A",X"C9",X"CD",X"BC",X"19",X"C0",X"FD",X"66",X"21",X"FD",X"6E",X"23",X"CD",
		X"F2",X"19",X"FE",X"FF",X"C8",X"B7",X"C9",X"FD",X"7E",X"16",X"B7",X"20",X"1A",X"3E",X"0C",X"16",
		X"00",X"1E",X"00",X"CD",X"20",X"2C",X"FD",X"7E",X"0E",X"FD",X"E5",X"FD",X"21",X"2B",X"4A",X"21",
		X"49",X"25",X"CD",X"61",X"1A",X"FD",X"E1",X"FD",X"7E",X"16",X"3C",X"FD",X"77",X"16",X"FE",X"10",
		X"28",X"10",X"FE",X"08",X"C0",X"FD",X"34",X"17",X"FD",X"34",X"17",X"FD",X"34",X"1B",X"FD",X"34",
		X"1B",X"C9",X"FD",X"36",X"17",X"00",X"FD",X"36",X"1B",X"00",X"3E",X"0C",X"CD",X"8E",X"2C",X"C3",
		X"AD",X"12",X"3E",X"15",X"FF",X"21",X"A1",X"4B",X"06",X"0F",X"CF",X"3E",X"3E",X"32",X"A2",X"4B",
		X"3C",X"32",X"A7",X"4B",X"3E",X"15",X"32",X"A4",X"4B",X"32",X"A9",X"4B",X"FD",X"7E",X"21",X"C6",
		X"F8",X"32",X"A3",X"4B",X"C6",X"10",X"32",X"A8",X"4B",X"FD",X"7E",X"23",X"D6",X"10",X"FE",X"10",
		X"30",X"02",X"3E",X"10",X"32",X"A5",X"4B",X"32",X"AA",X"4B",X"AF",X"32",X"A1",X"4B",X"32",X"A6",
		X"4B",X"FD",X"7E",X"0E",X"CD",X"E0",X"19",X"7C",X"32",X"8A",X"4B",X"32",X"8F",X"4B",X"32",X"94",
		X"4B",X"32",X"99",X"4B",X"32",X"9E",X"4B",X"7D",X"32",X"8C",X"4B",X"32",X"91",X"4B",X"32",X"96",
		X"4B",X"32",X"9B",X"4B",X"32",X"A0",X"4B",X"3E",X"18",X"32",X"9F",X"4B",X"3E",X"9F",X"32",X"8B",
		X"4B",X"32",X"90",X"4B",X"32",X"95",X"4B",X"32",X"9A",X"4B",X"21",X"55",X"25",X"11",X"14",X"4A",
		X"01",X"1A",X"00",X"ED",X"B0",X"3E",X"23",X"06",X"02",X"FF",X"FD",X"21",X"15",X"4A",X"DD",X"21",
		X"88",X"4B",X"06",X"04",X"C5",X"FD",X"7E",X"03",X"FD",X"B6",X"04",X"CA",X"4F",X"19",X"FD",X"7E",
		X"00",X"B7",X"28",X"05",X"FD",X"35",X"00",X"20",X"1E",X"FD",X"36",X"00",X"03",X"FD",X"6E",X"01",
		X"FD",X"66",X"02",X"7E",X"B7",X"20",X"06",X"01",X"08",X"00",X"ED",X"42",X"7E",X"23",X"FD",X"75",
		X"01",X"FD",X"74",X"02",X"DD",X"77",X"01",X"FD",X"6E",X"03",X"FD",X"66",X"04",X"7E",X"FE",X"80",
		X"20",X"16",X"FD",X"36",X"03",X"00",X"FD",X"36",X"04",X"00",X"3A",X"14",X"4A",X"3C",X"32",X"14",
		X"4A",X"FE",X"04",X"CA",X"95",X"19",X"18",X"37",X"4F",X"23",X"46",X"23",X"FD",X"75",X"03",X"FD",
		X"74",X"04",X"DD",X"66",X"02",X"DD",X"6E",X"04",X"CD",X"83",X"3D",X"7D",X"FE",X"10",X"30",X"04",
		X"2E",X"10",X"18",X"06",X"FE",X"FC",X"38",X"02",X"2E",X"FC",X"7C",X"FE",X"1C",X"30",X"04",X"26",
		X"1C",X"18",X"06",X"FE",X"F4",X"38",X"02",X"26",X"F4",X"DD",X"74",X"02",X"DD",X"75",X"04",X"DD",
		X"36",X"00",X"00",X"01",X"05",X"00",X"FD",X"09",X"DD",X"09",X"C1",X"05",X"C2",X"C4",X"18",X"FD",
		X"7E",X"00",X"B7",X"C2",X"B5",X"18",X"FD",X"7E",X"01",X"B7",X"28",X"06",X"FD",X"35",X"01",X"C3",
		X"B5",X"18",X"FD",X"6E",X"02",X"FD",X"66",X"03",X"7E",X"B7",X"20",X"03",X"FD",X"34",X"00",X"DD",
		X"77",X"01",X"23",X"7E",X"FD",X"77",X"01",X"23",X"FD",X"75",X"02",X"FD",X"74",X"03",X"DD",X"36",
		X"00",X"00",X"C3",X"B5",X"18",X"3E",X"23",X"06",X"10",X"FF",X"18",X"05",X"3E",X"23",X"06",X"40",
		X"FF",X"3E",X"47",X"06",X"20",X"FF",X"FD",X"21",X"14",X"4A",X"FD",X"6E",X"26",X"FD",X"66",X"27",
		X"3E",X"60",X"BE",X"20",X"04",X"FD",X"7E",X"29",X"77",X"3E",X"60",X"FF",X"FD",X"7E",X"21",X"E6",
		X"0F",X"C0",X"FD",X"7E",X"23",X"E6",X"0F",X"FE",X"08",X"C9",X"E6",X"0F",X"CD",X"F7",X"3D",X"21",
		X"9D",X"26",X"16",X"00",X"5F",X"19",X"7E",X"C9",X"21",X"4E",X"81",X"16",X"00",X"5F",X"19",X"C9",
		X"21",X"59",X"26",X"CD",X"E1",X"3D",X"D5",X"C1",X"FD",X"66",X"01",X"FD",X"6E",X"03",X"CD",X"83",
		X"3D",X"C9",X"E5",X"FD",X"7E",X"0E",X"21",X"61",X"26",X"CD",X"E1",X"3D",X"D5",X"C1",X"E1",X"CD",
		X"83",X"3D",X"CD",X"9E",X"0F",X"C9",X"FD",X"6E",X"0C",X"FD",X"66",X"0D",X"29",X"F5",X"11",X"00",
		X"00",X"ED",X"5A",X"FD",X"75",X"0C",X"FD",X"74",X"0D",X"F1",X"C9",X"FD",X"7E",X"0E",X"CD",X"E1",
		X"3D",X"EB",X"4E",X"23",X"46",X"23",X"5E",X"23",X"56",X"23",X"E5",X"FD",X"66",X"21",X"FD",X"6E",
		X"23",X"E5",X"CD",X"83",X"3D",X"FD",X"74",X"01",X"FD",X"75",X"03",X"E1",X"E5",X"D5",X"C1",X"CD",
		X"83",X"3D",X"FD",X"74",X"05",X"FD",X"75",X"07",X"D1",X"E1",X"3E",X"03",X"FD",X"BE",X"09",X"C0",
		X"4E",X"23",X"46",X"EB",X"CD",X"83",X"3D",X"FD",X"74",X"18",X"FD",X"75",X"1A",X"C9",X"FD",X"7E",
		X"0E",X"5F",X"87",X"83",X"16",X"00",X"5F",X"19",X"7E",X"23",X"FD",X"77",X"00",X"3C",X"FD",X"77",
		X"04",X"3A",X"1C",X"4A",X"FE",X"02",X"C8",X"7E",X"23",X"FD",X"77",X"20",X"3E",X"03",X"FD",X"BE",
		X"09",X"C0",X"7E",X"FD",X"77",X"17",X"C9",X"FD",X"7E",X"0A",X"21",X"69",X"26",X"CD",X"E1",X"3D",
		X"FD",X"73",X"0C",X"FD",X"72",X"0D",X"C9",X"FD",X"7E",X"0A",X"16",X"00",X"5F",X"21",X"AB",X"1A",
		X"19",X"FD",X"7E",X"10",X"E6",X"80",X"B6",X"FD",X"77",X"10",X"C9",X"0A",X"0A",X"0A",X"08",X"08",
		X"06",X"06",X"FD",X"7E",X"10",X"CB",X"BF",X"B7",X"28",X"04",X"FD",X"35",X"10",X"C9",X"CD",X"97",
		X"1A",X"21",X"7D",X"26",X"FD",X"7E",X"0E",X"CD",X"E1",X"3D",X"FD",X"CB",X"10",X"7E",X"20",X"17",
		X"7A",X"FD",X"BE",X"00",X"28",X"17",X"FD",X"CB",X"10",X"BE",X"FD",X"34",X"00",X"FD",X"34",X"00",
		X"FD",X"34",X"04",X"FD",X"34",X"04",X"C9",X"7B",X"FD",X"BE",X"00",X"28",X"E9",X"FD",X"CB",X"10",
		X"FE",X"FD",X"35",X"00",X"FD",X"35",X"00",X"FD",X"35",X"04",X"FD",X"35",X"04",X"C9",X"3A",X"01",
		X"48",X"CB",X"7F",X"28",X"17",X"21",X"00",X"50",X"3A",X"01",X"48",X"CB",X"6F",X"28",X"0A",X"3A",
		X"1B",X"48",X"CB",X"47",X"20",X"03",X"21",X"40",X"50",X"7E",X"2F",X"C9",X"C1",X"3A",X"42",X"4A",
		X"B7",X"28",X"10",X"3D",X"32",X"42",X"4A",X"28",X"0A",X"2A",X"40",X"4A",X"7E",X"FD",X"77",X"0F",
		X"C3",X"24",X"13",X"2A",X"40",X"4A",X"23",X"23",X"7E",X"FE",X"F0",X"28",X"0A",X"FE",X"F1",X"28",
		X"0C",X"CD",X"53",X"1B",X"C3",X"24",X"13",X"22",X"40",X"4A",X"C3",X"C2",X"12",X"22",X"40",X"4A",
		X"C3",X"29",X"16",X"22",X"40",X"4A",X"23",X"7E",X"32",X"42",X"4A",X"2B",X"7E",X"FD",X"77",X"0F",
		X"C9",X"3A",X"20",X"48",X"B7",X"C8",X"F5",X"CD",X"BB",X"1B",X"F1",X"CB",X"4F",X"C4",X"20",X"1D",
		X"C9",X"DD",X"21",X"58",X"4A",X"06",X"03",X"DD",X"7E",X"09",X"FE",X"04",X"30",X"24",X"FD",X"7E",
		X"21",X"C6",X"04",X"57",X"D6",X"08",X"5F",X"DD",X"7E",X"01",X"BA",X"30",X"15",X"BB",X"38",X"12",
		X"FD",X"7E",X"23",X"C6",X"04",X"57",X"D6",X"08",X"5F",X"DD",X"7E",X"03",X"BA",X"30",X"03",X"BB",
		X"30",X"08",X"11",X"30",X"00",X"DD",X"19",X"10",X"CE",X"C9",X"CD",X"6C",X"17",X"FD",X"E5",X"DD",
		X"E5",X"FD",X"E1",X"CD",X"84",X"24",X"FD",X"E1",X"DD",X"E1",X"C9",X"CD",X"E1",X"1C",X"C2",X"95",
		X"1C",X"CD",X"BA",X"1C",X"FE",X"FF",X"C8",X"E6",X"F0",X"C8",X"FE",X"70",X"D0",X"FD",X"E5",X"1A",
		X"FE",X"60",X"20",X"1D",X"E5",X"D5",X"3E",X"0D",X"CD",X"8E",X"2C",X"3A",X"01",X"48",X"F6",X"0A",
		X"32",X"01",X"48",X"CD",X"2B",X"1C",X"3E",X"06",X"01",X"28",X"86",X"FF",X"FD",X"7E",X"29",X"D1",
		X"E1",X"4F",X"E6",X"F0",X"FE",X"50",X"20",X"0B",X"FD",X"7E",X"09",X"FE",X"04",X"28",X"04",X"FD",
		X"36",X"09",X"02",X"79",X"E6",X"0F",X"12",X"CD",X"02",X"8D",X"FD",X"E1",X"3A",X"DB",X"49",X"3C",
		X"32",X"DB",X"49",X"3A",X"E0",X"49",X"3D",X"32",X"E0",X"49",X"28",X"05",X"FE",X"08",X"28",X"13",
		X"C9",X"3A",X"01",X"48",X"CB",X"4F",X"CB",X"CF",X"32",X"01",X"48",X"FD",X"36",X"0A",X"02",X"CD",
		X"87",X"1A",X"C9",X"3A",X"DA",X"49",X"CB",X"4F",X"C0",X"CB",X"4F",X"32",X"DA",X"49",X"3A",X"01",
		X"48",X"CB",X"67",X"CB",X"E7",X"32",X"01",X"48",X"3E",X"0D",X"16",X"00",X"1E",X"00",X"CD",X"20",
		X"2C",X"3A",X"01",X"48",X"CB",X"7F",X"20",X"05",X"21",X"57",X"48",X"18",X"1F",X"ED",X"5F",X"5F",
		X"16",X"00",X"21",X"30",X"48",X"19",X"B7",X"11",X"02",X"49",X"E5",X"ED",X"52",X"E1",X"38",X"03",
		X"21",X"30",X"48",X"7E",X"E6",X"F0",X"28",X"1A",X"FE",X"50",X"30",X"16",X"7E",X"FD",X"77",X"29",
		X"36",X"60",X"FD",X"75",X"26",X"FD",X"74",X"27",X"21",X"5A",X"02",X"FD",X"75",X"24",X"FD",X"74",
		X"25",X"C9",X"23",X"18",X"D1",X"21",X"10",X"1D",X"CD",X"E4",X"1C",X"C0",X"21",X"B2",X"1C",X"CD",
		X"BD",X"1C",X"47",X"FE",X"FF",X"C8",X"E6",X"F0",X"FE",X"90",X"D8",X"EB",X"CD",X"4A",X"17",X"C3",
		X"6C",X"17",X"00",X"F8",X"10",X"08",X"00",X"18",X"00",X"08",X"21",X"85",X"26",X"FD",X"7E",X"0E",
		X"CD",X"E1",X"3D",X"FD",X"7E",X"21",X"E6",X"F0",X"67",X"FD",X"7E",X"23",X"E6",X"F0",X"6F",X"D5",
		X"C1",X"CD",X"83",X"3D",X"E5",X"CD",X"BC",X"3D",X"D1",X"EB",X"D5",X"CD",X"9E",X"0F",X"D1",X"EB",
		X"C9",X"21",X"04",X"1D",X"FD",X"7E",X"0E",X"16",X"00",X"5F",X"87",X"83",X"5F",X"19",X"FD",X"CB",
		X"0E",X"46",X"FD",X"7E",X"21",X"20",X"03",X"FD",X"7E",X"23",X"E6",X"0F",X"BE",X"C8",X"23",X"BE",
		X"C8",X"23",X"BE",X"C9",X"05",X"06",X"07",X"01",X"02",X"03",X"09",X"0A",X"0B",X"0D",X"0E",X"0F",
		X"01",X"02",X"03",X"05",X"06",X"07",X"0D",X"0E",X"0F",X"09",X"0A",X"0B",X"FF",X"FF",X"FF",X"FF",
		X"3A",X"01",X"48",X"CB",X"4F",X"C0",X"C3",X"71",X"1B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"31",X"70",X"4E",X"21",X"56",X"4A",X"06",X"92",X"CF",X"21",X"A9",X"28",X"CD",X"84",X"24",X"FE",
		X"00",X"28",X"02",X"3E",X"01",X"CD",X"E1",X"3D",X"EB",X"46",X"23",X"FD",X"21",X"58",X"4A",X"C5",
		X"5E",X"23",X"56",X"23",X"E5",X"EB",X"FD",X"E5",X"D1",X"01",X"0D",X"00",X"ED",X"B0",X"21",X"80",
		X"00",X"FD",X"75",X"17",X"FD",X"74",X"18",X"11",X"30",X"00",X"FD",X"19",X"E1",X"C1",X"10",X"DF",
		X"3A",X"E3",X"49",X"B7",X"20",X"20",X"21",X"FA",X"28",X"CD",X"84",X"24",X"CD",X"E1",X"3D",X"EB",
		X"46",X"23",X"FD",X"21",X"24",X"48",X"5E",X"23",X"56",X"23",X"FD",X"73",X"00",X"FD",X"72",X"01",
		X"FD",X"23",X"FD",X"23",X"10",X"F0",X"AF",X"32",X"57",X"4A",X"3E",X"30",X"FF",X"3E",X"23",X"06",
		X"01",X"FF",X"FD",X"21",X"58",X"4A",X"DD",X"21",X"A1",X"4B",X"21",X"3E",X"28",X"CD",X"84",X"24",
		X"16",X"00",X"5F",X"19",X"46",X"AF",X"32",X"56",X"4A",X"C5",X"3A",X"01",X"48",X"E6",X"06",X"28",
		X"08",X"FD",X"7E",X"09",X"FE",X"04",X"DA",X"BF",X"1F",X"DD",X"E5",X"FD",X"7E",X"09",X"DF",X"EF",
		X"1D",X"9B",X"21",X"B4",X"21",X"6E",X"24",X"A4",X"20",X"07",X"21",X"D8",X"1F",X"2B",X"20",X"FD",
		X"7E",X"08",X"21",X"F8",X"1D",X"F7",X"18",X"0A",X"2C",X"21",X"2C",X"21",X"2C",X"21",X"2C",X"21",
		X"2C",X"21",X"FD",X"7E",X"08",X"FE",X"02",X"28",X"04",X"FE",X"03",X"20",X"54",X"FD",X"6E",X"17",
		X"FD",X"66",X"18",X"7D",X"B4",X"20",X"43",X"FD",X"7E",X"01",X"67",X"E6",X"0F",X"20",X"42",X"FD",
		X"7E",X"03",X"6F",X"E6",X"0F",X"FE",X"08",X"20",X"38",X"CD",X"C4",X"3F",X"38",X"33",X"21",X"60",
		X"27",X"CD",X"84",X"24",X"16",X"00",X"5F",X"19",X"FD",X"7E",X"19",X"3C",X"FD",X"77",X"19",X"BE",
		X"38",X"1F",X"AF",X"FD",X"77",X"19",X"21",X"6C",X"27",X"CD",X"84",X"24",X"CD",X"E1",X"3D",X"EB",
		X"3A",X"01",X"48",X"CB",X"7F",X"20",X"03",X"21",X"90",X"00",X"2B",X"FD",X"75",X"17",X"FD",X"74",
		X"18",X"3A",X"1D",X"4A",X"FE",X"04",X"C2",X"02",X"1F",X"3A",X"20",X"48",X"CB",X"5F",X"CA",X"02",
		X"1F",X"CD",X"7D",X"1E",X"D2",X"02",X"1F",X"21",X"5F",X"28",X"C3",X"7E",X"1F",X"3A",X"2C",X"4A",
		X"FD",X"BE",X"01",X"20",X"17",X"3A",X"2E",X"4A",X"C6",X"14",X"30",X"02",X"3E",X"FF",X"FD",X"BE",
		X"03",X"38",X"6D",X"C6",X"D8",X"FD",X"BE",X"03",X"30",X"66",X"18",X"49",X"3A",X"2E",X"4A",X"FD",
		X"BE",X"03",X"20",X"17",X"3A",X"2C",X"4A",X"C6",X"14",X"30",X"02",X"3E",X"FF",X"FD",X"BE",X"01",
		X"38",X"4E",X"C6",X"D8",X"FD",X"BE",X"01",X"30",X"47",X"18",X"2A",X"3A",X"2C",X"4A",X"C6",X"08",
		X"30",X"02",X"3E",X"FF",X"FD",X"BE",X"01",X"38",X"37",X"C6",X"F0",X"FD",X"BE",X"01",X"30",X"30",
		X"3A",X"2E",X"4A",X"C6",X"08",X"30",X"02",X"3E",X"FF",X"FD",X"BE",X"03",X"38",X"22",X"C6",X"F0",
		X"FD",X"BE",X"03",X"30",X"1B",X"3E",X"11",X"16",X"00",X"1E",X"00",X"CD",X"20",X"2C",X"FD",X"36",
		X"09",X"05",X"FD",X"36",X"0C",X"08",X"FD",X"36",X"00",X"34",X"FD",X"36",X"02",X"49",X"37",X"C9",
		X"A7",X"C9",X"FD",X"7E",X"14",X"B7",X"28",X"20",X"FD",X"35",X"14",X"C2",X"81",X"1F",X"FD",X"6E",
		X"15",X"FD",X"66",X"16",X"E5",X"CD",X"68",X"0F",X"E1",X"DD",X"E5",X"DD",X"21",X"77",X"89",X"1E",
		X"01",X"CD",X"50",X"89",X"DD",X"E1",X"18",X"59",X"3A",X"1C",X"4A",X"FE",X"03",X"20",X"52",X"3A",
		X"22",X"4A",X"EE",X"02",X"FD",X"BE",X"0A",X"20",X"48",X"3A",X"35",X"4A",X"C6",X"02",X"FD",X"BE",
		X"01",X"38",X"3E",X"D6",X"04",X"FD",X"BE",X"01",X"30",X"37",X"3A",X"37",X"4A",X"C6",X"02",X"FD",
		X"BE",X"03",X"38",X"2D",X"D6",X"04",X"FD",X"BE",X"03",X"30",X"26",X"FD",X"66",X"01",X"FD",X"6E",
		X"03",X"CD",X"9E",X"0F",X"CD",X"F4",X"0F",X"FD",X"75",X"15",X"FD",X"74",X"16",X"FD",X"36",X"14",
		X"40",X"3E",X"CC",X"1E",X"15",X"01",X"02",X"02",X"CD",X"1E",X"3D",X"21",X"59",X"28",X"CD",X"04",
		X"3E",X"DD",X"E1",X"FD",X"E5",X"E1",X"DD",X"E5",X"D1",X"13",X"01",X"04",X"00",X"ED",X"B0",X"FD",
		X"7E",X"09",X"FE",X"06",X"20",X"04",X"DD",X"36",X"01",X"00",X"DD",X"36",X"00",X"00",X"3A",X"01",
		X"48",X"CB",X"7F",X"28",X"1A",X"3A",X"56",X"4A",X"21",X"24",X"48",X"CD",X"E1",X"3D",X"3A",X"DC",
		X"49",X"47",X"1A",X"B8",X"20",X"09",X"13",X"1A",X"FD",X"77",X"08",X"13",X"72",X"2B",X"73",X"3A",
		X"56",X"4A",X"3C",X"32",X"56",X"4A",X"01",X"30",X"00",X"FD",X"09",X"01",X"05",X"00",X"DD",X"09",
		X"C1",X"05",X"C2",X"C9",X"1D",X"C3",X"AD",X"1D",X"FD",X"6E",X"0B",X"FD",X"66",X"0C",X"2B",X"FD",
		X"75",X"0B",X"FD",X"74",X"0C",X"7D",X"B4",X"C2",X"81",X"1F",X"CD",X"62",X"20",X"FD",X"36",X"09",
		X"07",X"3A",X"01",X"48",X"CB",X"7F",X"20",X"19",X"3A",X"57",X"4A",X"F5",X"21",X"84",X"27",X"CD",
		X"E1",X"3D",X"F1",X"3C",X"32",X"57",X"4A",X"FD",X"73",X"1A",X"FD",X"72",X"1B",X"AF",X"FD",X"77",
		X"1C",X"21",X"8B",X"20",X"FD",X"75",X"0D",X"FD",X"74",X"0E",X"3E",X"11",X"CD",X"8E",X"2C",X"3E",
		X"06",X"16",X"00",X"1E",X"00",X"CD",X"20",X"2C",X"C3",X"81",X"1F",X"FD",X"7E",X"0C",X"B7",X"28",
		X"06",X"FD",X"35",X"0C",X"C3",X"81",X"1F",X"FD",X"36",X"0C",X"0A",X"FD",X"6E",X"0D",X"FD",X"66",
		X"0E",X"7E",X"FE",X"FF",X"28",X"12",X"23",X"5E",X"23",X"FD",X"75",X"0D",X"FD",X"74",X"0E",X"FD",
		X"77",X"00",X"FD",X"73",X"02",X"C3",X"81",X"1F",X"CD",X"62",X"20",X"FD",X"36",X"09",X"00",X"C3",
		X"81",X"1F",X"FD",X"7E",X"08",X"F5",X"21",X"A9",X"28",X"CD",X"84",X"24",X"FE",X"00",X"28",X"02",
		X"3E",X"01",X"CD",X"E1",X"3D",X"EB",X"23",X"3A",X"56",X"4A",X"CD",X"E1",X"3D",X"EB",X"FD",X"E5",
		X"D1",X"01",X"0B",X"00",X"ED",X"B0",X"F1",X"FD",X"77",X"08",X"C9",X"29",X"08",X"2F",X"5C",X"30",
		X"5B",X"29",X"08",X"2F",X"5B",X"30",X"5C",X"29",X"5B",X"2F",X"08",X"30",X"5C",X"29",X"5B",X"2F",
		X"08",X"30",X"5C",X"FF",X"CD",X"AA",X"20",X"C3",X"81",X"1F",X"FD",X"7E",X"0C",X"B7",X"20",X"08",
		X"FD",X"36",X"00",X"25",X"FD",X"36",X"02",X"4F",X"3C",X"FD",X"77",X"0C",X"FE",X"40",X"C0",X"FD",
		X"36",X"09",X"06",X"FD",X"36",X"00",X"00",X"3A",X"56",X"4A",X"CB",X"27",X"CB",X"27",X"21",X"FB",
		X"20",X"16",X"00",X"5F",X"19",X"3E",X"02",X"01",X"C0",X"00",X"F5",X"5E",X"23",X"56",X"23",X"1A",
		X"FE",X"06",X"20",X"0C",X"E5",X"13",X"13",X"EB",X"5E",X"23",X"56",X"EB",X"09",X"4D",X"44",X"E1",
		X"F1",X"3D",X"20",X"E6",X"FD",X"71",X"0B",X"FD",X"70",X"0C",X"C9",X"91",X"4A",X"C1",X"4A",X"61",
		X"4A",X"C1",X"4A",X"61",X"4A",X"91",X"4A",X"CD",X"0D",X"21",X"C3",X"81",X"1F",X"FD",X"35",X"0C",
		X"C0",X"FD",X"36",X"0C",X"08",X"FD",X"7E",X"00",X"3C",X"FD",X"77",X"00",X"FE",X"37",X"C0",X"FD",
		X"36",X"00",X"00",X"FD",X"36",X"0C",X"00",X"FD",X"36",X"09",X"04",X"C9",X"3E",X"01",X"FD",X"BE",
		X"09",X"28",X"06",X"21",X"A1",X"28",X"CD",X"AD",X"80",X"3A",X"01",X"48",X"CB",X"7F",X"CA",X"D7",
		X"22",X"FD",X"7E",X"01",X"E6",X"0F",X"C2",X"85",X"21",X"FD",X"7E",X"03",X"E6",X"0F",X"FE",X"08",
		X"C2",X"85",X"21",X"FD",X"7E",X"11",X"B7",X"CA",X"B6",X"22",X"3E",X"01",X"FD",X"BE",X"08",X"20",
		X"12",X"3A",X"8A",X"4B",X"FD",X"BE",X"01",X"CA",X"B6",X"22",X"3A",X"8C",X"4B",X"FD",X"BE",X"03",
		X"CA",X"B6",X"22",X"CD",X"8E",X"24",X"FD",X"7E",X"0A",X"CD",X"EB",X"3D",X"FD",X"A6",X"13",X"CA",
		X"B6",X"22",X"C3",X"00",X"80",X"FD",X"7E",X"0A",X"CD",X"EB",X"3D",X"F5",X"CD",X"9A",X"24",X"CD",
		X"5A",X"81",X"F1",X"A1",X"C2",X"00",X"80",X"CD",X"6E",X"24",X"C9",X"FD",X"7E",X"0B",X"B7",X"28",
		X"06",X"FD",X"35",X"0B",X"C3",X"EF",X"1D",X"FD",X"36",X"09",X"00",X"21",X"9D",X"28",X"CD",X"64",
		X"80",X"C3",X"EF",X"1D",X"FD",X"7E",X"12",X"B7",X"20",X"0E",X"FD",X"34",X"12",X"3E",X"01",X"FD",
		X"77",X"04",X"CD",X"81",X"80",X"CD",X"91",X"80",X"21",X"A1",X"28",X"CD",X"AD",X"80",X"FD",X"7E",
		X"01",X"E6",X"0F",X"20",X"5C",X"FD",X"7E",X"03",X"E6",X"0F",X"FE",X"08",X"20",X"53",X"CD",X"8E",
		X"24",X"FD",X"7E",X"08",X"FE",X"02",X"28",X"5D",X"3E",X"0A",X"FD",X"CB",X"0A",X"46",X"28",X"02",
		X"3E",X"05",X"FD",X"A6",X"13",X"28",X"2D",X"FD",X"77",X"13",X"FD",X"36",X"09",X"00",X"21",X"4A",
		X"28",X"CD",X"70",X"80",X"3A",X"01",X"48",X"CB",X"7F",X"20",X"06",X"CD",X"D7",X"22",X"C3",X"02",
		X"1E",X"3E",X"01",X"FD",X"BE",X"08",X"20",X"06",X"CD",X"14",X"23",X"C3",X"02",X"1E",X"CD",X"B9",
		X"22",X"C3",X"02",X"1E",X"FD",X"7E",X"0A",X"EE",X"02",X"CD",X"EB",X"3D",X"FD",X"A6",X"13",X"28",
		X"06",X"CD",X"00",X"80",X"C3",X"02",X"1E",X"FD",X"7E",X"0A",X"CD",X"EB",X"3D",X"FD",X"A6",X"13",
		X"CA",X"02",X"1E",X"18",X"B5",X"21",X"AE",X"22",X"FD",X"7E",X"0A",X"CD",X"E1",X"3D",X"06",X"05",
		X"0E",X"0F",X"FD",X"66",X"01",X"FD",X"6E",X"03",X"C5",X"D5",X"E5",X"CD",X"9E",X"0F",X"FE",X"FF",
		X"28",X"09",X"47",X"E6",X"F0",X"28",X"06",X"FE",X"80",X"28",X"02",X"AF",X"47",X"78",X"E6",X"0F",
		X"21",X"4E",X"81",X"16",X"00",X"5F",X"19",X"7E",X"E1",X"D1",X"C1",X"A1",X"4F",X"FD",X"CB",X"0A",
		X"46",X"20",X"0B",X"7D",X"FE",X"18",X"28",X"18",X"FE",X"F8",X"28",X"14",X"18",X"09",X"7C",X"FE",
		X"20",X"28",X"0D",X"FE",X"F0",X"28",X"09",X"C5",X"D5",X"C1",X"CD",X"83",X"3D",X"C1",X"10",X"B8",
		X"FD",X"7E",X"0A",X"59",X"CD",X"EB",X"3D",X"A3",X"C2",X"FA",X"21",X"C3",X"E8",X"21",X"00",X"F0",
		X"10",X"00",X"00",X"10",X"F0",X"00",X"CD",X"8E",X"24",X"3A",X"01",X"48",X"CB",X"7F",X"CA",X"D7",
		X"22",X"3A",X"1D",X"4A",X"FE",X"01",X"CA",X"14",X"23",X"FD",X"7E",X"08",X"DF",X"14",X"23",X"DE",
		X"23",X"53",X"24",X"8D",X"23",X"53",X"24",X"FD",X"7E",X"1C",X"B7",X"28",X"08",X"FD",X"35",X"1C",
		X"28",X"03",X"C3",X"00",X"80",X"FD",X"6E",X"1A",X"FD",X"66",X"1B",X"23",X"23",X"FD",X"75",X"1A",
		X"FD",X"74",X"1B",X"7E",X"E6",X"F0",X"28",X"13",X"FE",X"F0",X"28",X"03",X"C3",X"6E",X"24",X"23",
		X"7E",X"FD",X"77",X"08",X"23",X"FD",X"75",X"1A",X"FD",X"74",X"1B",X"7E",X"23",X"46",X"FD",X"70",
		X"1C",X"C3",X"61",X"23",X"CD",X"E9",X"80",X"1E",X"00",X"FD",X"CB",X"0A",X"46",X"20",X"02",X"1E",
		X"01",X"CB",X"4F",X"28",X"04",X"7B",X"C6",X"02",X"5F",X"7B",X"CD",X"EB",X"3D",X"FD",X"A6",X"13",
		X"20",X"1A",X"7B",X"EE",X"02",X"CD",X"EB",X"3D",X"FD",X"A6",X"13",X"20",X"0F",X"FD",X"7E",X"0A",
		X"CD",X"EB",X"3D",X"FD",X"A6",X"13",X"20",X"04",X"CD",X"6E",X"24",X"C9",X"F5",X"CD",X"E9",X"80",
		X"E6",X"0F",X"21",X"8D",X"28",X"16",X"00",X"5F",X"19",X"7E",X"FD",X"77",X"11",X"F1",X"CD",X"F7",
		X"3D",X"FD",X"BE",X"0A",X"CA",X"00",X"80",X"FD",X"77",X"0B",X"21",X"60",X"28",X"FD",X"7E",X"0A",
		X"CD",X"E1",X"3D",X"EB",X"FD",X"7E",X"0B",X"FD",X"77",X"0A",X"16",X"00",X"5F",X"19",X"7E",X"FD",
		X"77",X"00",X"FD",X"36",X"09",X"01",X"FD",X"36",X"0B",X"08",X"C3",X"00",X"80",X"CD",X"59",X"24",
		X"16",X"40",X"3A",X"22",X"4A",X"CB",X"47",X"20",X"20",X"CB",X"4F",X"20",X"08",X"7D",X"92",X"30",
		X"0C",X"3E",X"18",X"30",X"08",X"7D",X"82",X"30",X"04",X"3E",X"F8",X"18",X"00",X"6F",X"7C",X"26",
		X"D0",X"FE",X"80",X"38",X"02",X"26",X"40",X"18",X"1C",X"CB",X"4F",X"20",X"08",X"7C",X"82",X"30",
		X"0A",X"3E",X"F0",X"18",X"06",X"7C",X"92",X"30",X"02",X"3E",X"20",X"67",X"7D",X"2E",X"40",X"FE",
		X"80",X"30",X"02",X"2E",X"D0",X"FD",X"74",X"0F",X"FD",X"75",X"10",X"C3",X"C0",X"87",X"CD",X"59",
		X"24",X"FD",X"7E",X"0A",X"CD",X"EB",X"3D",X"47",X"FD",X"CB",X"0A",X"46",X"20",X"24",X"FD",X"7E",
		X"01",X"FD",X"BE",X"0F",X"20",X"07",X"78",X"FD",X"A6",X"13",X"C2",X"4C",X"23",X"06",X"02",X"FD",
		X"7E",X"01",X"FD",X"BE",X"0F",X"38",X"02",X"06",X"08",X"78",X"FD",X"A6",X"13",X"C2",X"4C",X"23",
		X"18",X"22",X"FD",X"7E",X"03",X"FD",X"BE",X"10",X"20",X"07",X"78",X"FD",X"A6",X"13",X"C2",X"4C",
		X"23",X"06",X"01",X"FD",X"7E",X"03",X"FD",X"BE",X"10",X"30",X"02",X"06",X"04",X"78",X"FD",X"A6",
		X"13",X"C2",X"4C",X"23",X"78",X"CD",X"F7",X"3D",X"EE",X"02",X"CD",X"EB",X"3D",X"FD",X"A6",X"13",
		X"C2",X"4C",X"23",X"FD",X"7E",X"0A",X"CD",X"EB",X"3D",X"FD",X"A6",X"13",X"C2",X"4C",X"23",X"CD",
		X"6E",X"24",X"C9",X"CD",X"59",X"24",X"C3",X"C0",X"87",X"3A",X"35",X"4A",X"E6",X"F0",X"FD",X"77",
		X"0F",X"67",X"3A",X"37",X"4A",X"E6",X"F0",X"C6",X"08",X"FD",X"77",X"10",X"6F",X"C9",X"FD",X"7E",
		X"09",X"FE",X"01",X"20",X"06",X"21",X"9D",X"28",X"CD",X"64",X"80",X"FD",X"36",X"09",X"02",X"FD",
		X"36",X"12",X"00",X"C9",X"3A",X"E7",X"49",X"FE",X"0C",X"D8",X"D6",X"0C",X"18",X"F9",X"3E",X"0F",
		X"F5",X"CD",X"FD",X"80",X"F1",X"A1",X"FD",X"77",X"13",X"C9",X"3A",X"56",X"4A",X"21",X"78",X"28",
		X"CD",X"E1",X"3D",X"EB",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"02",X"10",X"01",X"20",X"04",X"40",X"F0",X"00",X"04",X"10",X"01",X"10",X"04",X"10",X"08",X"18",
		X"F1",X"00",X"01",X"28",X"02",X"40",X"F0",X"00",X"02",X"10",X"08",X"60",X"04",X"40",X"08",X"40",
		X"04",X"50",X"01",X"08",X"F1",X"00",X"01",X"28",X"02",X"30",X"F0",X"00",X"01",X"30",X"01",X"40",
		X"04",X"50",X"08",X"10",X"F0",X"00",X"02",X"10",X"01",X"20",X"02",X"30",X"F0",X"00",X"08",X"10",
		X"04",X"90",X"08",X"10",X"02",X"10",X"08",X"10",X"02",X"10",X"08",X"40",X"02",X"20",X"01",X"50",
		X"02",X"60",X"08",X"10",X"02",X"10",X"01",X"20",X"72",X"73",X"A7",X"A8",X"32",X"33",X"27",X"28",
		X"00",X"FC",X"04",X"00",X"00",X"04",X"FC",X"00",X"5A",X"5A",X"5A",X"5A",X"5A",X"5A",X"5A",X"5A",
		X"5A",X"5A",X"00",X"FF",X"01",X"00",X"00",X"01",X"FF",X"00",X"00",X"FE",X"02",X"00",X"00",X"02",
		X"FE",X"00",X"01",X"02",X"03",X"04",X"00",X"01",X"0B",X"15",X"00",X"00",X"19",X"00",X"00",X"15",
		X"00",X"00",X"19",X"00",X"00",X"00",X"00",X"6E",X"25",X"80",X"25",X"00",X"77",X"25",X"BD",X"25",
		X"00",X"6E",X"25",X"FA",X"25",X"00",X"77",X"25",X"1F",X"26",X"00",X"00",X"44",X"26",X"3B",X"BC",
		X"BD",X"FC",X"7B",X"7C",X"3D",X"3C",X"00",X"3B",X"3C",X"3D",X"7C",X"7B",X"FC",X"BD",X"BC",X"00",
		X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",
		X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",
		X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",
		X"00",X"01",X"FF",X"01",X"00",X"01",X"FF",X"01",X"00",X"01",X"00",X"01",X"80",X"01",X"FE",X"01",
		X"FE",X"01",X"FE",X"01",X"FE",X"01",X"FE",X"01",X"FE",X"01",X"FE",X"01",X"FE",X"01",X"FE",X"01",
		X"FE",X"01",X"FE",X"01",X"FE",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"00",X"01",X"00",X"01",
		X"00",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"01",X"01",
		X"01",X"00",X"01",X"01",X"01",X"00",X"01",X"00",X"01",X"80",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",
		X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"FF",X"00",
		X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"80",X"02",
		X"FF",X"02",X"FF",X"02",X"FF",X"02",X"FF",X"02",X"FF",X"02",X"FF",X"02",X"FF",X"01",X"00",X"01",
		X"00",X"01",X"00",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"80",X"39",X"06",X"38",X"06",X"37",X"06",X"38",X"06",X"39",X"06",X"38",X"06",
		X"37",X"06",X"38",X"06",X"39",X"06",X"38",X"06",X"00",X"00",X"08",X"F8",X"00",X"00",X"F8",X"08",
		X"00",X"00",X"F0",X"10",X"00",X"00",X"10",X"F0",X"00",X"00",X"00",X"22",X"22",X"55",X"55",X"D6",
		X"D6",X"EE",X"EE",X"FE",X"FE",X"FF",X"FF",X"80",X"80",X"88",X"88",X"AA",X"AA",X"41",X"43",X"85",
		X"87",X"01",X"03",X"05",X"07",X"00",X"F8",X"10",X"08",X"00",X"18",X"00",X"08",X"95",X"26",X"99",
		X"26",X"95",X"26",X"99",X"26",X"F8",X"00",X"08",X"00",X"00",X"F8",X"00",X"08",X"00",X"03",X"01",
		X"02",X"04",X"AA",X"26",X"B6",X"26",X"C2",X"26",X"CE",X"26",X"00",X"00",X"00",X"C9",X"E3",X"00",
		X"01",X"1D",X"00",X"49",X"63",X"00",X"8B",X"A4",X"00",X"00",X"00",X"00",X"CB",X"E4",X"00",X"05",
		X"1E",X"00",X"41",X"5D",X"00",X"89",X"A3",X"00",X"00",X"00",X"00",X"09",X"23",X"00",X"0B",X"24",
		X"00",X"85",X"9E",X"00",X"4B",X"64",X"00",X"00",X"00",X"00",X"E2",X"26",X"E8",X"26",X"EE",X"26",
		X"F4",X"26",X"00",X"F8",X"00",X"08",X"00",X"F0",X"08",X"00",X"F8",X"00",X"10",X"00",X"00",X"08",
		X"00",X"F8",X"00",X"10",X"F8",X"00",X"08",X"00",X"F0",X"00",X"41",X"5D",X"71",X"85",X"9E",X"A6",
		X"01",X"1D",X"31",X"05",X"1E",X"26",X"0A",X"27",X"16",X"27",X"4F",X"60",X"00",X"93",X"A2",X"00",
		X"0F",X"20",X"00",X"13",X"22",X"00",X"4D",X"5F",X"00",X"91",X"A1",X"00",X"0D",X"1F",X"00",X"11",
		X"21",X"00",X"05",X"78",X"9F",X"98",X"06",X"88",X"9F",X"98",X"00",X"00",X"02",X"02",X"AA",X"AA",
		X"03",X"04",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"1E",X"80",X"9E",X"98",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"04",X"03",X"02",X"03",X"01",X"02",X"01",X"02",X"01",X"03",X"01",X"01",X"B0",X"00",X"80",X"00",
		X"40",X"00",X"60",X"00",X"20",X"00",X"20",X"00",X"40",X"00",X"40",X"00",X"20",X"00",X"40",X"00",
		X"30",X"00",X"30",X"00",X"88",X"27",X"8E",X"27",X"DE",X"27",X"F0",X"00",X"01",X"10",X"00",X"FF",
		X"01",X"10",X"02",X"10",X"03",X"40",X"00",X"10",X"03",X"10",X"02",X"10",X"E0",X"00",X"01",X"10",
		X"02",X"10",X"F0",X"02",X"01",X"40",X"02",X"30",X"03",X"10",X"00",X"10",X"03",X"40",X"02",X"20",
		X"03",X"10",X"02",X"10",X"03",X"10",X"02",X"20",X"01",X"10",X"02",X"10",X"01",X"10",X"00",X"10",
		X"01",X"40",X"00",X"20",X"03",X"30",X"02",X"10",X"01",X"30",X"00",X"10",X"01",X"10",X"00",X"60",
		X"03",X"40",X"F0",X"00",X"02",X"10",X"01",X"40",X"02",X"90",X"03",X"20",X"00",X"10",X"01",X"30",
		X"F0",X"00",X"01",X"10",X"00",X"60",X"03",X"40",X"02",X"10",X"03",X"60",X"02",X"10",X"03",X"20",
		X"02",X"30",X"03",X"10",X"02",X"10",X"01",X"70",X"00",X"10",X"03",X"10",X"E0",X"00",X"02",X"10",
		X"03",X"30",X"00",X"70",X"01",X"40",X"02",X"10",X"01",X"30",X"02",X"20",X"01",X"10",X"02",X"20",
		X"03",X"20",X"1A",X"28",X"23",X"28",X"2C",X"28",X"35",X"28",X"EC",X"AD",X"AC",X"2A",X"2C",X"2D",
		X"6C",X"6A",X"00",X"AC",X"2A",X"2C",X"2D",X"6C",X"6A",X"EC",X"AD",X"00",X"2C",X"2D",X"6C",X"6A",
		X"EC",X"AD",X"AC",X"2A",X"00",X"6C",X"6A",X"EC",X"AD",X"AC",X"2A",X"2C",X"2D",X"00",X"02",X"03",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"06",X"06",X"06",X"06",X"06",X"06",
		X"06",X"06",X"06",X"06",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"68",X"28",X"6C",X"28",X"70",X"28",X"74",X"28",X"00",X"EC",X"2A",X"6C",X"EC",X"00",X"AC",X"2D",
		X"6A",X"AC",X"00",X"2C",X"6C",X"AD",X"2C",X"00",X"7E",X"28",X"83",X"28",X"88",X"28",X"02",X"88",
		X"4A",X"B8",X"4A",X"02",X"58",X"4A",X"B8",X"4A",X"02",X"58",X"4A",X"88",X"4A",X"10",X"20",X"30",
		X"10",X"50",X"40",X"10",X"30",X"20",X"10",X"40",X"50",X"10",X"20",X"10",X"30",X"6A",X"AD",X"2A",
		X"2D",X"6A",X"6B",X"AD",X"AE",X"2A",X"2B",X"2D",X"2E",X"AD",X"28",X"B2",X"28",X"02",X"B9",X"28",
		X"C6",X"28",X"03",X"D3",X"28",X"E0",X"28",X"ED",X"28",X"AD",X"E0",X"5B",X"B8",X"06",X"06",X"FF",
		X"FF",X"02",X"06",X"01",X"3C",X"00",X"AD",X"A0",X"5C",X"18",X"06",X"06",X"FF",X"FF",X"03",X"06",
		X"01",X"B4",X"00",X"6A",X"F0",X"5B",X"F8",X"06",X"06",X"FF",X"FF",X"03",X"06",X"00",X"3C",X"00",
		X"AD",X"A0",X"5C",X"18",X"06",X"06",X"FF",X"FF",X"01",X"06",X"01",X"B4",X"00",X"AD",X"20",X"5D",
		X"F8",X"06",X"06",X"FF",X"FF",X"02",X"06",X"01",X"2D",X"01",X"12",X"29",X"17",X"29",X"1E",X"29",
		X"25",X"29",X"2C",X"29",X"33",X"29",X"3A",X"29",X"41",X"29",X"48",X"29",X"4F",X"29",X"56",X"29",
		X"5D",X"29",X"02",X"64",X"29",X"75",X"29",X"03",X"86",X"29",X"9B",X"29",X"AE",X"29",X"03",X"C1",
		X"29",X"D2",X"29",X"E3",X"29",X"03",X"F6",X"29",X"0D",X"2A",X"1E",X"2A",X"03",X"2F",X"2A",X"46",
		X"2A",X"57",X"2A",X"03",X"68",X"2A",X"7F",X"2A",X"90",X"2A",X"03",X"A1",X"2A",X"B8",X"2A",X"C9",
		X"2A",X"03",X"DA",X"2A",X"F1",X"2A",X"02",X"2B",X"03",X"13",X"2B",X"2A",X"2B",X"3B",X"2B",X"03",
		X"4C",X"2B",X"65",X"2B",X"78",X"2B",X"03",X"8F",X"2B",X"A6",X"2B",X"BD",X"2B",X"03",X"D4",X"2B",
		X"ED",X"2B",X"04",X"2C",X"00",X"01",X"0A",X"02",X"14",X"02",X"1E",X"01",X"28",X"02",X"32",X"03",
		X"37",X"02",X"46",X"02",X"FF",X"00",X"03",X"0A",X"01",X"14",X"00",X"1E",X"01",X"28",X"03",X"32",
		X"00",X"3C",X"01",X"46",X"01",X"FF",X"00",X"03",X"0A",X"02",X"14",X"03",X"1E",X"00",X"28",X"02",
		X"30",X"01",X"32",X"01",X"3C",X"03",X"46",X"01",X"50",X"01",X"FF",X"00",X"00",X"0A",X"01",X"14",
		X"00",X"1E",X"02",X"28",X"01",X"30",X"02",X"3C",X"03",X"46",X"02",X"50",X"02",X"FF",X"00",X"02",
		X"0A",X"03",X"14",X"01",X"1E",X"01",X"28",X"03",X"32",X"01",X"3C",X"00",X"46",X"01",X"50",X"01",
		X"FF",X"00",X"01",X"0A",X"02",X"14",X"00",X"1E",X"01",X"32",X"03",X"3C",X"01",X"32",X"03",X"32",
		X"03",X"FF",X"00",X"02",X"14",X"03",X"1E",X"02",X"28",X"01",X"32",X"02",X"3C",X"03",X"46",X"02",
		X"50",X"02",X"FF",X"00",X"00",X"0A",X"01",X"14",X"01",X"1E",X"00",X"28",X"02",X"32",X"01",X"3C",
		X"00",X"41",X"01",X"50",X"01",X"FF",X"00",X"00",X"08",X"01",X"0A",X"02",X"14",X"03",X"1E",X"02",
		X"28",X"00",X"32",X"01",X"3C",X"02",X"46",X"01",X"50",X"02",X"5A",X"02",X"FF",X"00",X"01",X"0A",
		X"01",X"1E",X"03",X"28",X"02",X"3C",X"01",X"46",X"01",X"50",X"03",X"5A",X"01",X"FF",X"00",X"02",
		X"0A",X"03",X"14",X"02",X"28",X"01",X"32",X"03",X"3C",X"01",X"4B",X"00",X"50",X"01",X"FF",X"00",
		X"01",X"08",X"01",X"0A",X"02",X"14",X"03",X"1E",X"02",X"28",X"00",X"32",X"01",X"3C",X"02",X"46",
		X"02",X"50",X"03",X"5A",X"02",X"FF",X"00",X"01",X"0A",X"01",X"1E",X"03",X"28",X"02",X"3C",X"01",
		X"46",X"01",X"55",X"00",X"5A",X"01",X"FF",X"00",X"02",X"0A",X"03",X"14",X"02",X"28",X"00",X"32",
		X"01",X"3C",X"03",X"46",X"01",X"50",X"01",X"FF",X"00",X"01",X"08",X"01",X"0A",X"02",X"14",X"03",
		X"1E",X"02",X"28",X"00",X"32",X"01",X"3C",X"02",X"46",X"02",X"50",X"03",X"5A",X"02",X"FF",X"00",
		X"01",X"0A",X"01",X"1E",X"04",X"28",X"02",X"3C",X"01",X"46",X"01",X"50",X"02",X"5A",X"01",X"FF",
		X"00",X"02",X"0A",X"03",X"14",X"02",X"28",X"00",X"32",X"01",X"3C",X"01",X"46",X"04",X"50",X"01",
		X"FF",X"00",X"04",X"08",X"04",X"0A",X"02",X"14",X"04",X"1E",X"02",X"28",X"00",X"32",X"01",X"3C",
		X"02",X"46",X"02",X"50",X"01",X"5A",X"02",X"FF",X"00",X"01",X"0A",X"01",X"1E",X"03",X"28",X"02",
		X"3C",X"01",X"46",X"01",X"50",X"02",X"5A",X"01",X"FF",X"00",X"02",X"0A",X"03",X"14",X"02",X"28",
		X"04",X"32",X"01",X"3C",X"01",X"46",X"01",X"50",X"04",X"FF",X"00",X"04",X"08",X"01",X"0A",X"02",
		X"14",X"03",X"1E",X"02",X"28",X"04",X"32",X"01",X"3C",X"02",X"46",X"02",X"50",X"01",X"5A",X"02",
		X"FF",X"00",X"01",X"0A",X"01",X"1E",X"03",X"28",X"02",X"3C",X"01",X"46",X"01",X"50",X"02",X"5A",
		X"01",X"FF",X"00",X"02",X"0A",X"03",X"14",X"02",X"28",X"00",X"32",X"01",X"3C",X"01",X"46",X"01",
		X"50",X"04",X"FF",X"00",X"04",X"08",X"04",X"0A",X"02",X"14",X"03",X"1E",X"02",X"28",X"00",X"32",
		X"01",X"3C",X"02",X"46",X"02",X"50",X"01",X"5A",X"02",X"FF",X"00",X"01",X"0A",X"01",X"1E",X"04",
		X"28",X"02",X"3C",X"01",X"46",X"01",X"50",X"02",X"5A",X"01",X"FF",X"00",X"02",X"0A",X"03",X"14",
		X"02",X"28",X"00",X"32",X"04",X"3C",X"01",X"46",X"01",X"50",X"04",X"FF",X"00",X"04",X"08",X"04",
		X"0A",X"02",X"14",X"03",X"1E",X"02",X"28",X"00",X"2D",X"04",X"32",X"01",X"3C",X"02",X"46",X"02",
		X"50",X"01",X"5A",X"02",X"FF",X"00",X"04",X"0A",X"01",X"1E",X"04",X"23",X"00",X"28",X"02",X"3C",
		X"01",X"46",X"01",X"50",X"02",X"5A",X"01",X"FF",X"00",X"02",X"0A",X"03",X"14",X"02",X"1E",X"00",
		X"23",X"04",X"28",X"04",X"2D",X"00",X"32",X"04",X"3C",X"01",X"46",X"01",X"50",X"04",X"FF",X"00",
		X"04",X"08",X"04",X"0A",X"02",X"14",X"03",X"1E",X"02",X"28",X"00",X"32",X"01",X"3C",X"02",X"46",
		X"02",X"50",X"01",X"5A",X"02",X"FF",X"00",X"01",X"0A",X"01",X"14",X"00",X"19",X"04",X"1E",X"04",
		X"23",X"00",X"28",X"02",X"3C",X"01",X"46",X"01",X"50",X"02",X"5A",X"01",X"FF",X"00",X"02",X"0A",
		X"03",X"14",X"02",X"1E",X"00",X"23",X"00",X"28",X"04",X"32",X"04",X"37",X"00",X"3C",X"01",X"46",
		X"01",X"50",X"04",X"FF",X"00",X"04",X"08",X"04",X"0A",X"02",X"14",X"03",X"1E",X"02",X"28",X"00",
		X"32",X"01",X"3C",X"02",X"41",X"00",X"46",X"02",X"50",X"01",X"5A",X"02",X"FF",X"00",X"01",X"0A",
		X"01",X"0F",X"00",X"14",X"04",X"1E",X"04",X"23",X"00",X"28",X"02",X"3C",X"01",X"46",X"01",X"50",
		X"02",X"5A",X"01",X"FF",X"00",X"02",X"0A",X"03",X"14",X"02",X"28",X"00",X"32",X"04",X"3C",X"01",
		X"41",X"00",X"46",X"01",X"50",X"04",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"08",X"28",X"08",X"47",X"3A",X"01",X"48",X"CB",X"7F",X"C8",X"78",X"DD",X"E5",X"FD",X"E5",
		X"CD",X"EE",X"2C",X"CD",X"D9",X"2C",X"DD",X"7E",X"00",X"E6",X"0F",X"D5",X"CD",X"C9",X"2C",X"D1",
		X"C5",X"E5",X"06",X"10",X"CD",X"58",X"2D",X"E1",X"C1",X"E5",X"23",X"DD",X"7E",X"01",X"83",X"77",
		X"23",X"DD",X"7E",X"02",X"82",X"77",X"23",X"FD",X"E5",X"E5",X"FD",X"E1",X"DD",X"7E",X"03",X"77",
		X"FD",X"77",X"03",X"23",X"DD",X"7E",X"04",X"77",X"FD",X"77",X"04",X"FD",X"E1",X"23",X"3E",X"01",
		X"77",X"E1",X"DD",X"7E",X"00",X"E6",X"40",X"F6",X"80",X"77",X"DD",X"CB",X"00",X"7E",X"20",X"09",
		X"C5",X"01",X"05",X"00",X"DD",X"09",X"C1",X"18",X"AD",X"FD",X"E1",X"DD",X"E1",X"C9",X"DD",X"E5",
		X"FD",X"E5",X"CD",X"EE",X"2C",X"CD",X"D9",X"2C",X"DD",X"7E",X"00",X"E6",X"0F",X"47",X"CB",X"20",
		X"CD",X"C9",X"2C",X"CB",X"66",X"C4",X"91",X"2E",X"C5",X"06",X"10",X"CD",X"58",X"2D",X"C1",X"11",
		X"00",X"80",X"CD",X"D7",X"2F",X"16",X"8F",X"CD",X"E2",X"2F",X"DD",X"CB",X"00",X"7E",X"20",X"C9",
		X"C5",X"01",X"05",X"00",X"DD",X"09",X"C1",X"18",X"CF",X"21",X"D6",X"2C",X"5F",X"16",X"00",X"19",
		X"5E",X"FD",X"E5",X"E1",X"19",X"C9",X"00",X"10",X"20",X"21",X"00",X"4C",X"B7",X"28",X"0B",X"D5",
		X"C5",X"11",X"30",X"00",X"47",X"19",X"10",X"FD",X"C1",X"D1",X"E5",X"FD",X"E1",X"C9",X"87",X"87",
		X"4F",X"06",X"00",X"DD",X"21",X"12",X"31",X"DD",X"09",X"DD",X"7E",X"00",X"DD",X"4E",X"01",X"DD",
		X"6E",X"02",X"DD",X"66",X"03",X"E5",X"DD",X"E1",X"C9",X"06",X"02",X"3E",X"00",X"C5",X"F5",X"CD",
		X"18",X"2D",X"F1",X"C1",X"3C",X"10",X"F6",X"C9",X"F5",X"CD",X"D9",X"2C",X"06",X"30",X"CD",X"58",
		X"2D",X"F1",X"CD",X"4D",X"2D",X"2E",X"03",X"06",X"00",X"16",X"8F",X"CD",X"E2",X"2F",X"11",X"00",
		X"80",X"CD",X"D7",X"2F",X"04",X"04",X"2D",X"20",X"F0",X"06",X"06",X"CD",X"DF",X"2F",X"2E",X"04",
		X"06",X"00",X"16",X"8F",X"CD",X"E2",X"2F",X"04",X"04",X"2D",X"20",X"F8",X"C9",X"21",X"10",X"31",
		X"D5",X"5F",X"16",X"00",X"19",X"D1",X"4E",X"C9",X"36",X"00",X"23",X"10",X"FB",X"C9",X"06",X"02",
		X"3E",X"00",X"FD",X"21",X"00",X"4C",X"F5",X"C5",X"CD",X"4D",X"2D",X"06",X"00",X"FD",X"CB",X"00",
		X"7E",X"C5",X"C4",X"88",X"2D",X"C1",X"11",X"10",X"00",X"FD",X"19",X"04",X"04",X"78",X"FE",X"06",
		X"20",X"EB",X"C1",X"F1",X"3C",X"10",X"DF",X"C9",X"FD",X"CB",X"00",X"6E",X"C2",X"2E",X"2F",X"FD",
		X"CB",X"00",X"5E",X"C2",X"3F",X"2F",X"FD",X"35",X"05",X"C0",X"FD",X"7E",X"02",X"FD",X"77",X"05",
		X"FD",X"CB",X"00",X"4E",X"28",X"08",X"FD",X"35",X"0D",X"C0",X"FD",X"CB",X"00",X"8E",X"FD",X"CB",
		X"00",X"46",X"28",X"0E",X"FD",X"35",X"0D",X"C0",X"FD",X"56",X"0F",X"CD",X"E2",X"2F",X"FD",X"CB",
		X"00",X"86",X"FD",X"6E",X"06",X"FD",X"66",X"07",X"7E",X"23",X"FD",X"75",X"06",X"FD",X"74",X"07",
		X"CB",X"7F",X"20",X"29",X"C5",X"47",X"E6",X"0F",X"87",X"4F",X"78",X"0F",X"0F",X"0F",X"0F",X"E6",
		X"07",X"FD",X"86",X"01",X"6F",X"26",X"00",X"29",X"29",X"29",X"E5",X"D1",X"19",X"19",X"11",X"F6",
		X"2F",X"06",X"00",X"19",X"09",X"C1",X"56",X"23",X"5E",X"CD",X"D7",X"2F",X"C9",X"F5",X"E6",X"8F",
		X"57",X"F1",X"D5",X"07",X"07",X"07",X"07",X"E6",X"07",X"21",X"18",X"2E",X"16",X"00",X"CB",X"27",
		X"5F",X"19",X"5E",X"23",X"56",X"EB",X"D1",X"E9",X"28",X"2E",X"3C",X"2E",X"50",X"2E",X"59",X"2E",
		X"64",X"2E",X"A0",X"2E",X"B6",X"2E",X"A3",X"2F",X"7A",X"E6",X"07",X"CB",X"62",X"28",X"02",X"ED",
		X"44",X"57",X"FD",X"7E",X"02",X"82",X"FD",X"77",X"02",X"C3",X"C2",X"2D",X"7A",X"E6",X"07",X"CB",
		X"62",X"28",X"02",X"ED",X"44",X"57",X"FD",X"7E",X"01",X"82",X"FD",X"77",X"01",X"C3",X"C2",X"2D",
		X"FD",X"72",X"0F",X"CD",X"E2",X"2F",X"C3",X"C2",X"2D",X"7A",X"E6",X"0F",X"FD",X"77",X"0D",X"FD",
		X"CB",X"00",X"CE",X"C9",X"7A",X"FE",X"8F",X"28",X"1E",X"FD",X"CB",X"00",X"E6",X"C5",X"06",X"06",
		X"CD",X"E2",X"2F",X"FD",X"6E",X"06",X"FD",X"66",X"07",X"7E",X"57",X"23",X"FD",X"75",X"06",X"FD",
		X"74",X"07",X"CD",X"DF",X"2F",X"C1",X"C9",X"FD",X"CB",X"00",X"A6",X"CD",X"91",X"2E",X"C3",X"C2",
		X"2D",X"C5",X"06",X"06",X"16",X"8F",X"CD",X"E2",X"2F",X"16",X"80",X"CD",X"DF",X"2F",X"C1",X"C9",
		X"7A",X"E6",X"0F",X"FD",X"77",X"0D",X"FD",X"CB",X"00",X"C6",X"16",X"8F",X"CD",X"E2",X"2F",X"11",
		X"00",X"80",X"CD",X"D7",X"2F",X"C9",X"FD",X"6E",X"06",X"FD",X"66",X"07",X"2B",X"7E",X"FE",X"E0",
		X"28",X"3C",X"7A",X"E6",X"0F",X"21",X"B8",X"30",X"3D",X"87",X"5F",X"16",X"00",X"19",X"5E",X"23",
		X"56",X"EB",X"FD",X"7E",X"02",X"FD",X"77",X"0D",X"FD",X"77",X"0E",X"FD",X"75",X"0B",X"FD",X"74",
		X"0C",X"FD",X"6E",X"06",X"FD",X"66",X"07",X"7E",X"23",X"FD",X"75",X"06",X"FD",X"74",X"07",X"FD",
		X"CB",X"00",X"EE",X"CD",X"D4",X"2D",X"FD",X"6E",X"0B",X"FD",X"66",X"0C",X"18",X"71",X"23",X"7E",
		X"FD",X"77",X"0D",X"FD",X"77",X"0E",X"23",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"FD",X"75",X"0B",
		X"FD",X"74",X"0C",X"5F",X"16",X"00",X"19",X"7E",X"23",X"FD",X"CB",X"00",X"DE",X"FD",X"75",X"06",
		X"FD",X"74",X"07",X"CD",X"D4",X"2D",X"FD",X"6E",X"0B",X"FD",X"66",X"0C",X"18",X"41",X"FD",X"35",
		X"05",X"C0",X"FD",X"35",X"0E",X"FD",X"6E",X"0B",X"FD",X"66",X"0C",X"20",X"32",X"18",X"53",X"FD",
		X"35",X"05",X"C8",X"FD",X"35",X"0E",X"FD",X"6E",X"0B",X"FD",X"66",X"0C",X"20",X"21",X"FD",X"7E",
		X"0D",X"FD",X"77",X"0E",X"FD",X"6E",X"06",X"FD",X"66",X"07",X"7E",X"23",X"FD",X"75",X"06",X"FD",
		X"74",X"07",X"FE",X"E0",X"28",X"2C",X"CD",X"D4",X"2D",X"FD",X"6E",X"09",X"FD",X"66",X"0A",X"7E",
		X"F5",X"23",X"FD",X"75",X"0B",X"FD",X"74",X"0C",X"07",X"07",X"07",X"07",X"E6",X"0F",X"FD",X"77",
		X"05",X"FD",X"7E",X"0F",X"E6",X"0F",X"57",X"F1",X"E6",X"0F",X"82",X"F6",X"80",X"57",X"CD",X"E2",
		X"2F",X"C9",X"FD",X"CB",X"00",X"9E",X"FD",X"CB",X"00",X"AE",X"FD",X"7E",X"02",X"FD",X"77",X"05",
		X"C3",X"C2",X"2D",X"FD",X"CB",X"00",X"BE",X"FD",X"CB",X"00",X"66",X"FD",X"CB",X"00",X"A6",X"C4",
		X"91",X"2E",X"16",X"8F",X"CD",X"E2",X"2F",X"11",X"00",X"80",X"CD",X"D7",X"2F",X"FD",X"CB",X"00",
		X"76",X"C8",X"FD",X"36",X"00",X"C0",X"FD",X"6E",X"03",X"FD",X"66",X"04",X"FD",X"75",X"06",X"FD",
		X"74",X"07",X"FD",X"36",X"05",X"01",X"C9",X"CD",X"E9",X"2F",X"7B",X"CD",X"F3",X"2F",X"C9",X"57",
		X"18",X"07",X"C5",X"04",X"CD",X"E9",X"2F",X"C1",X"C9",X"78",X"07",X"07",X"07",X"07",X"B2",X"CD",
		X"F3",X"2F",X"C9",X"ED",X"79",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"88",X"3F",X"8F",X"3B",X"89",X"38",X"86",X"35",X"86",X"32",X"8A",X"2F",X"8E",X"2C",X"86",X"2A",
		X"80",X"28",X"8C",X"25",X"8A",X"23",X"8A",X"21",X"8C",X"1F",X"8F",X"1D",X"84",X"1C",X"8B",X"1A",
		X"83",X"19",X"8D",X"17",X"87",X"16",X"83",X"15",X"80",X"14",X"8E",X"12",X"8D",X"11",X"8D",X"10",
		X"8E",X"0F",X"80",X"0F",X"82",X"0E",X"86",X"0D",X"8A",X"0C",X"8E",X"0B",X"84",X"0B",X"8A",X"0A",
		X"80",X"0A",X"87",X"09",X"8F",X"08",X"87",X"08",X"8F",X"07",X"88",X"07",X"81",X"07",X"8B",X"06",
		X"85",X"06",X"8F",X"05",X"8A",X"05",X"85",X"05",X"80",X"05",X"8B",X"04",X"87",X"04",X"83",X"04",
		X"8F",X"03",X"8C",X"03",X"89",X"03",X"86",X"03",X"83",X"03",X"80",X"03",X"8D",X"02",X"8B",X"02",
		X"88",X"02",X"86",X"02",X"83",X"02",X"82",X"02",X"8F",X"01",X"8E",X"01",X"8C",X"01",X"8B",X"01",
		X"8A",X"01",X"88",X"01",X"87",X"01",X"86",X"01",X"84",X"01",X"82",X"01",X"81",X"01",X"80",X"01",
		X"8F",X"00",X"8E",X"00",X"8D",X"00",X"FF",X"FF",X"C8",X"30",X"D1",X"30",X"DA",X"30",X"E3",X"30",
		X"EC",X"30",X"F5",X"30",X"FE",X"30",X"07",X"31",X"80",X"82",X"80",X"82",X"80",X"82",X"80",X"82",
		X"80",X"40",X"42",X"40",X"42",X"40",X"42",X"40",X"42",X"40",X"20",X"22",X"20",X"22",X"20",X"22",
		X"20",X"22",X"20",X"10",X"12",X"10",X"12",X"10",X"12",X"10",X"12",X"10",X"80",X"81",X"82",X"83",
		X"84",X"85",X"86",X"87",X"88",X"40",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"48",X"20",X"21",
		X"22",X"23",X"24",X"25",X"26",X"27",X"28",X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"18",
		X"01",X"02",X"01",X"02",X"5A",X"31",X"00",X"01",X"79",X"32",X"00",X"01",X"A5",X"32",X"00",X"01",
		X"D1",X"32",X"01",X"02",X"FD",X"32",X"00",X"01",X"0D",X"33",X"00",X"01",X"1E",X"33",X"01",X"02",
		X"3A",X"33",X"00",X"01",X"71",X"33",X"00",X"01",X"8B",X"33",X"00",X"01",X"AF",X"33",X"00",X"01",
		X"E0",X"33",X"01",X"02",X"27",X"34",X"00",X"01",X"4B",X"34",X"00",X"01",X"8D",X"34",X"00",X"01",
		X"A7",X"34",X"01",X"02",X"EE",X"34",X"00",X"01",X"01",X"35",X"40",X"00",X"05",X"64",X"31",X"C1",
		X"00",X"05",X"EF",X"31",X"A7",X"D4",X"E3",X"34",X"E3",X"2B",X"E3",X"32",X"E3",X"33",X"D2",X"E3",
		X"34",X"D2",X"E3",X"37",X"E3",X"39",X"E3",X"32",X"E3",X"37",X"E3",X"39",X"D4",X"D4",X"E1",X"44",
		X"E3",X"42",X"E3",X"44",X"E2",X"42",X"E3",X"3B",X"E3",X"42",X"E3",X"3A",X"E4",X"39",X"E4",X"37",
		X"E3",X"34",X"E3",X"32",X"D4",X"E3",X"39",X"E3",X"34",X"E3",X"37",X"E3",X"38",X"D2",X"E3",X"39",
		X"D2",X"E3",X"3B",X"E3",X"42",X"E3",X"3B",X"E3",X"42",X"E3",X"43",X"D4",X"D4",X"E1",X"44",X"E3",
		X"42",X"E3",X"44",X"E2",X"42",X"E3",X"3B",X"E3",X"42",X"E3",X"3A",X"E4",X"39",X"E4",X"37",X"E3",
		X"34",X"E3",X"32",X"D4",X"E2",X"42",X"D2",X"E3",X"3B",X"D4",X"E2",X"39",X"D2",X"E3",X"37",X"D2",
		X"E3",X"2B",X"E3",X"32",X"E3",X"33",X"E2",X"34",X"E1",X"44",X"E3",X"42",X"E3",X"44",X"E2",X"42",
		X"E3",X"3B",X"E3",X"42",X"E3",X"3A",X"E4",X"39",X"E4",X"37",X"E3",X"34",X"E3",X"32",X"FF",X"A6",
		X"E6",X"24",X"E7",X"24",X"E7",X"1B",X"D2",X"E7",X"1B",X"E6",X"22",X"E6",X"24",X"E7",X"24",X"E7",
		X"1B",X"D2",X"E7",X"1B",X"E6",X"22",X"E6",X"24",X"E7",X"24",X"E7",X"1B",X"D2",X"E7",X"1B",X"E6",
		X"22",X"E6",X"24",X"E7",X"24",X"E7",X"1B",X"D2",X"E7",X"1B",X"E6",X"22",X"E6",X"29",X"E7",X"29",
		X"E7",X"24",X"D2",X"E7",X"24",X"E6",X"27",X"E6",X"29",X"E7",X"29",X"E7",X"24",X"D2",X"E7",X"24",
		X"E6",X"27",X"E6",X"24",X"E7",X"24",X"E7",X"1B",X"D2",X"E7",X"1B",X"E6",X"22",X"E6",X"24",X"E7",
		X"24",X"E7",X"1B",X"D2",X"E7",X"1B",X"E6",X"22",X"E6",X"2B",X"E7",X"2B",X"E7",X"26",X"D2",X"E7",
		X"26",X"E7",X"2B",X"E7",X"2A",X"E6",X"29",X"E7",X"29",X"E7",X"24",X"D2",X"E7",X"24",X"E7",X"29",
		X"E7",X"27",X"E6",X"24",X"E7",X"24",X"E7",X"1B",X"D2",X"E7",X"1B",X"E6",X"22",X"E6",X"24",X"E7",
		X"24",X"E7",X"1B",X"D2",X"E7",X"1B",X"E6",X"22",X"FF",X"01",X"00",X"01",X"83",X"32",X"82",X"00",
		X"01",X"94",X"32",X"AA",X"40",X"A9",X"40",X"A6",X"40",X"A3",X"40",X"A4",X"40",X"A7",X"40",X"A9",
		X"40",X"AB",X"40",X"FF",X"AA",X"37",X"A9",X"37",X"A6",X"37",X"A3",X"37",X"A4",X"37",X"A7",X"37",
		X"A9",X"37",X"AB",X"37",X"FF",X"01",X"00",X"01",X"AF",X"32",X"82",X"00",X"01",X"C0",X"32",X"AA",
		X"44",X"A9",X"44",X"A6",X"44",X"A3",X"44",X"A4",X"44",X"A7",X"44",X"A9",X"44",X"AB",X"44",X"FF",
		X"AA",X"40",X"A9",X"40",X"A6",X"40",X"A3",X"40",X"A4",X"40",X"A7",X"40",X"A9",X"40",X"AB",X"40",
		X"FF",X"01",X"00",X"01",X"DB",X"32",X"82",X"00",X"01",X"EC",X"32",X"AA",X"47",X"A9",X"47",X"A6",
		X"47",X"A3",X"47",X"A4",X"47",X"A7",X"47",X"A9",X"47",X"AB",X"47",X"FF",X"AA",X"44",X"A9",X"44",
		X"A6",X"44",X"A3",X"44",X"A4",X"44",X"A7",X"44",X"A9",X"44",X"AB",X"44",X"FF",X"82",X"00",X"03",
		X"02",X"33",X"C0",X"87",X"7B",X"C6",X"87",X"78",X"CA",X"87",X"77",X"CF",X"FF",X"C1",X"00",X"02",
		X"12",X"33",X"A3",X"68",X"64",X"67",X"63",X"66",X"62",X"65",X"61",X"64",X"60",X"FF",X"82",X"00",
		X"04",X"23",X"33",X"A4",X"E0",X"04",X"24",X"20",X"23",X"26",X"28",X"25",X"29",X"26",X"2A",X"27",
		X"2B",X"28",X"30",X"29",X"31",X"2A",X"32",X"2B",X"E0",X"FF",X"82",X"00",X"01",X"3F",X"33",X"A3",
		X"20",X"35",X"21",X"36",X"22",X"37",X"23",X"38",X"24",X"39",X"25",X"3A",X"26",X"3B",X"27",X"40",
		X"28",X"41",X"29",X"42",X"2A",X"43",X"2B",X"44",X"2B",X"44",X"2A",X"43",X"29",X"42",X"28",X"41",
		X"27",X"40",X"26",X"3B",X"25",X"3A",X"24",X"39",X"23",X"38",X"22",X"37",X"21",X"36",X"20",X"35",
		X"FF",X"80",X"00",X"01",X"76",X"33",X"A4",X"4B",X"43",X"4B",X"43",X"D2",X"57",X"55",X"57",X"55",
		X"D2",X"54",X"51",X"54",X"51",X"D2",X"52",X"48",X"52",X"48",X"FF",X"81",X"00",X"05",X"90",X"33",
		X"A2",X"57",X"B5",X"D2",X"50",X"B5",X"D4",X"57",X"B5",X"D2",X"50",X"B5",X"D4",X"57",X"B5",X"D2",
		X"50",X"B5",X"D4",X"57",X"B5",X"D2",X"50",X"B5",X"D4",X"57",X"B5",X"D2",X"50",X"B5",X"FF",X"40",
		X"00",X"02",X"B9",X"33",X"C1",X"00",X"05",X"C2",X"33",X"A5",X"58",X"50",X"55",X"49",X"54",X"48",
		X"53",X"FF",X"A6",X"45",X"46",X"47",X"48",X"49",X"4A",X"4B",X"50",X"51",X"52",X"53",X"54",X"55",
		X"56",X"57",X"58",X"59",X"5A",X"5B",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"BF",X"FF",
		X"01",X"00",X"02",X"EA",X"33",X"82",X"00",X"06",X"04",X"34",X"A8",X"DF",X"65",X"6B",X"64",X"6A",
		X"63",X"69",X"62",X"68",X"61",X"67",X"60",X"66",X"5B",X"65",X"5A",X"64",X"59",X"63",X"58",X"62",
		X"57",X"61",X"56",X"FF",X"C0",X"86",X"1B",X"C2",X"84",X"1B",X"AF",X"C4",X"84",X"1A",X"C6",X"84",
		X"20",X"CF",X"C0",X"86",X"1B",X"CF",X"C3",X"86",X"1B",X"CF",X"C6",X"86",X"1B",X"CF",X"C9",X"86",
		X"1B",X"CF",X"C9",X"86",X"1B",X"CF",X"FF",X"82",X"00",X"04",X"2C",X"34",X"C0",X"82",X"1B",X"CF",
		X"C0",X"82",X"C1",X"82",X"1B",X"CF",X"C3",X"82",X"1B",X"CF",X"C5",X"82",X"1B",X"CF",X"C7",X"82",
		X"1B",X"CF",X"C9",X"82",X"1B",X"CF",X"CB",X"82",X"1B",X"CF",X"FF",X"40",X"00",X"04",X"55",X"34",
		X"C1",X"00",X"04",X"71",X"34",X"A4",X"E0",X"0B",X"49",X"47",X"45",X"43",X"41",X"40",X"41",X"43",
		X"45",X"47",X"49",X"57",X"B5",X"50",X"B5",X"57",X"B5",X"50",X"B5",X"57",X"B5",X"50",X"B5",X"E0",
		X"FF",X"A4",X"E0",X"0B",X"49",X"47",X"45",X"43",X"41",X"40",X"41",X"43",X"45",X"47",X"49",X"50",
		X"B5",X"44",X"B5",X"50",X"B5",X"44",X"B5",X"50",X"B5",X"44",X"B5",X"E0",X"FF",X"81",X"00",X"02",
		X"92",X"34",X"A3",X"E0",X"04",X"40",X"31",X"32",X"36",X"45",X"49",X"52",X"45",X"55",X"55",X"48",
		X"48",X"53",X"46",X"50",X"49",X"E0",X"FF",X"01",X"00",X"02",X"B1",X"34",X"82",X"00",X"02",X"CF",
		X"34",X"A8",X"78",X"77",X"75",X"74",X"73",X"72",X"71",X"70",X"6B",X"6A",X"69",X"68",X"67",X"66",
		X"65",X"64",X"63",X"62",X"61",X"60",X"5B",X"5A",X"59",X"58",X"57",X"56",X"55",X"54",X"FF",X"A6",
		X"C0",X"85",X"20",X"CF",X"C2",X"85",X"20",X"CF",X"C6",X"87",X"75",X"74",X"73",X"72",X"71",X"70",
		X"6B",X"6A",X"69",X"68",X"67",X"66",X"65",X"64",X"63",X"62",X"61",X"60",X"CF",X"FF",X"82",X"00",
		X"06",X"F3",X"34",X"C0",X"87",X"70",X"C1",X"87",X"70",X"C3",X"87",X"70",X"C5",X"87",X"70",X"CF",
		X"FF",X"82",X"00",X"06",X"06",X"35",X"C0",X"86",X"1B",X"CF",X"C3",X"86",X"1B",X"CF",X"C6",X"86",
		X"1B",X"CF",X"C9",X"86",X"1B",X"CF",X"C9",X"86",X"1B",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"31",X"90",X"4F",X"18",X"05",X"31",X"90",X"4F",X"18",X"1C",X"CD",X"09",X"2D",X"3A",X"80",X"50",
		X"2F",X"32",X"1B",X"48",X"CD",X"54",X"39",X"CD",X"79",X"39",X"21",X"FF",X"3B",X"11",X"00",X"B8",
		X"01",X"80",X"00",X"ED",X"B0",X"EF",X"21",X"DF",X"38",X"CD",X"A8",X"3D",X"21",X"02",X"48",X"36",
		X"00",X"2B",X"7E",X"E6",X"80",X"77",X"F5",X"3E",X"10",X"FF",X"CD",X"B0",X"39",X"CD",X"E6",X"38",
		X"CD",X"54",X"39",X"F1",X"CB",X"7F",X"CA",X"4A",X"36",X"3A",X"06",X"48",X"B7",X"20",X"0C",X"3A",
		X"04",X"48",X"B7",X"20",X"06",X"AF",X"32",X"01",X"48",X"18",X"CB",X"CD",X"F2",X"39",X"CD",X"71",
		X"3A",X"CD",X"23",X"3A",X"DD",X"21",X"F1",X"3A",X"CD",X"B2",X"3C",X"3A",X"1B",X"48",X"E6",X"C0",
		X"07",X"07",X"21",X"1D",X"3B",X"CD",X"E1",X"3D",X"D5",X"DD",X"E1",X"CD",X"B2",X"3C",X"DD",X"21",
		X"07",X"3B",X"CD",X"B2",X"3C",X"21",X"49",X"42",X"DD",X"21",X"07",X"48",X"1E",X"0B",X"06",X"02",
		X"0E",X"00",X"CD",X"8A",X"3D",X"3E",X"23",X"06",X"01",X"FF",X"3A",X"06",X"48",X"B7",X"20",X"09",
		X"DD",X"21",X"C7",X"3A",X"CD",X"B2",X"3C",X"18",X"EC",X"FE",X"02",X"30",X"1C",X"DD",X"21",X"90",
		X"3A",X"CD",X"B2",X"3C",X"3A",X"04",X"48",X"B7",X"28",X"07",X"DD",X"21",X"D7",X"3A",X"CD",X"B2",
		X"3C",X"06",X"20",X"18",X"14",X"00",X"01",X"00",X"02",X"DD",X"21",X"90",X"3A",X"CD",X"B2",X"3C",
		X"DD",X"21",X"AB",X"3A",X"CD",X"B2",X"3C",X"06",X"60",X"3A",X"40",X"50",X"2F",X"A0",X"CA",X"C5",
		X"35",X"21",X"01",X"48",X"11",X"F6",X"35",X"CB",X"27",X"CB",X"27",X"30",X"05",X"CB",X"F6",X"11",
		X"F8",X"35",X"23",X"CB",X"FE",X"EB",X"3A",X"06",X"48",X"96",X"32",X"06",X"48",X"11",X"08",X"48",
		X"06",X"02",X"CD",X"64",X"3D",X"21",X"49",X"42",X"DD",X"21",X"07",X"48",X"1E",X"0B",X"06",X"02",
		X"0E",X"00",X"CD",X"8A",X"3D",X"3E",X"23",X"06",X"04",X"FF",X"3A",X"01",X"48",X"CB",X"7F",X"20",
		X"22",X"3A",X"02",X"48",X"CB",X"77",X"CB",X"F7",X"32",X"02",X"48",X"CD",X"E9",X"38",X"21",X"30",
		X"48",X"CD",X"00",X"03",X"79",X"32",X"E0",X"49",X"CD",X"28",X"83",X"21",X"01",X"48",X"36",X"00",
		X"23",X"36",X"00",X"21",X"0F",X"48",X"06",X"0C",X"CF",X"21",X"90",X"39",X"11",X"D4",X"49",X"01",
		X"20",X"00",X"ED",X"B0",X"21",X"90",X"39",X"11",X"F4",X"49",X"01",X"20",X"00",X"ED",X"B0",X"21",
		X"30",X"48",X"CD",X"00",X"03",X"79",X"32",X"E0",X"49",X"21",X"02",X"49",X"CD",X"00",X"03",X"79",
		X"32",X"00",X"4A",X"3A",X"1B",X"48",X"E6",X"30",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"C6",X"03",X"32",X"E6",X"49",X"32",X"06",X"4A",X"CD",X"B0",X"39",X"CD",X"54",X"39",X"3E",X"10",
		X"FF",X"CD",X"F2",X"39",X"CD",X"71",X"3A",X"3A",X"01",X"48",X"CB",X"7F",X"28",X"06",X"3E",X"00",
		X"01",X"D8",X"85",X"FF",X"3A",X"E6",X"49",X"47",X"CD",X"EF",X"3E",X"21",X"40",X"42",X"01",X"0C",
		X"01",X"3E",X"00",X"1E",X"0A",X"CD",X"31",X"3D",X"18",X"03",X"CD",X"DE",X"39",X"3A",X"E3",X"49",
		X"B7",X"28",X"0E",X"CD",X"E6",X"38",X"CD",X"15",X"39",X"3E",X"23",X"06",X"60",X"FF",X"CD",X"DE",
		X"39",X"CD",X"E9",X"38",X"DD",X"21",X"B0",X"3B",X"CD",X"B2",X"3C",X"DD",X"21",X"14",X"3B",X"CD",
		X"B2",X"3C",X"21",X"20",X"41",X"DD",X"21",X"E8",X"49",X"1E",X"0A",X"06",X"02",X"0E",X"FF",X"CD",
		X"8A",X"3D",X"CD",X"12",X"3F",X"3A",X"E3",X"49",X"B7",X"28",X"08",X"CD",X"5C",X"0D",X"CD",X"E9",
		X"0E",X"18",X"0B",X"CD",X"5C",X"0D",X"3E",X"23",X"06",X"40",X"FF",X"CD",X"57",X"0E",X"3E",X"23",
		X"06",X"20",X"FF",X"21",X"D8",X"38",X"CD",X"B0",X"3D",X"CD",X"E9",X"0E",X"3E",X"30",X"FF",X"3E",
		X"80",X"FF",X"F5",X"21",X"DF",X"38",X"CD",X"A8",X"3D",X"CD",X"09",X"2D",X"21",X"01",X"48",X"7E",
		X"E6",X"E0",X"77",X"23",X"7E",X"E6",X"80",X"77",X"F1",X"FE",X"10",X"CA",X"67",X"38",X"3E",X"23",
		X"06",X"20",X"FF",X"3A",X"01",X"48",X"CB",X"7F",X"20",X"0C",X"CD",X"DE",X"39",X"CD",X"E6",X"38",
		X"CD",X"73",X"8B",X"C3",X"56",X"35",X"3A",X"E1",X"49",X"B7",X"20",X"17",X"21",X"90",X"39",X"11",
		X"D4",X"49",X"01",X"11",X"00",X"ED",X"B0",X"21",X"30",X"48",X"CD",X"00",X"03",X"79",X"32",X"E0",
		X"49",X"18",X"04",X"21",X"E3",X"49",X"34",X"21",X"E6",X"49",X"3A",X"01",X"48",X"CB",X"77",X"20",
		X"18",X"35",X"C2",X"EA",X"36",X"CD",X"F5",X"38",X"3E",X"23",X"06",X"80",X"FF",X"CD",X"DE",X"39",
		X"CD",X"E6",X"38",X"CD",X"90",X"8A",X"C3",X"56",X"35",X"35",X"20",X"13",X"CD",X"F5",X"38",X"3E",
		X"23",X"06",X"80",X"FF",X"CD",X"DE",X"39",X"CD",X"E6",X"38",X"CD",X"90",X"8A",X"18",X"07",X"3A",
		X"06",X"4A",X"B7",X"CA",X"EA",X"36",X"3A",X"06",X"4A",X"B7",X"CA",X"56",X"35",X"3A",X"01",X"48",
		X"CB",X"6F",X"CB",X"EF",X"28",X"02",X"CB",X"AF",X"32",X"01",X"48",X"21",X"30",X"48",X"11",X"14",
		X"4A",X"01",X"D2",X"00",X"ED",X"B0",X"21",X"02",X"49",X"11",X"30",X"48",X"01",X"D2",X"00",X"ED",
		X"B0",X"21",X"14",X"4A",X"11",X"02",X"49",X"01",X"D2",X"00",X"ED",X"B0",X"21",X"D4",X"49",X"11",
		X"14",X"4A",X"01",X"20",X"00",X"ED",X"B0",X"21",X"F4",X"49",X"11",X"D4",X"49",X"01",X"20",X"00",
		X"ED",X"B0",X"21",X"14",X"4A",X"11",X"F4",X"49",X"01",X"20",X"00",X"ED",X"B0",X"21",X"24",X"48",
		X"11",X"14",X"4A",X"01",X"06",X"00",X"ED",X"B0",X"21",X"2A",X"48",X"11",X"24",X"48",X"01",X"06",
		X"00",X"ED",X"B0",X"21",X"14",X"4A",X"11",X"2A",X"48",X"01",X"06",X"00",X"ED",X"B0",X"21",X"14",
		X"4A",X"06",X"D2",X"CF",X"C3",X"B8",X"36",X"3E",X"0A",X"16",X"00",X"1E",X"00",X"CD",X"20",X"2C",
		X"3A",X"E1",X"49",X"B7",X"28",X"1A",X"3D",X"32",X"E1",X"49",X"CD",X"12",X"3F",X"21",X"8F",X"38",
		X"CD",X"04",X"3E",X"3E",X"23",X"06",X"03",X"FF",X"18",X"E6",X"00",X"00",X"00",X"00",X"05",X"00",
		X"3E",X"0A",X"CD",X"8E",X"2C",X"3E",X"23",X"06",X"20",X"FF",X"3A",X"01",X"48",X"CB",X"7F",X"CA",
		X"56",X"35",X"21",X"90",X"39",X"11",X"D4",X"49",X"01",X"11",X"00",X"ED",X"B0",X"21",X"D5",X"38",
		X"3A",X"E7",X"49",X"3C",X"FE",X"60",X"38",X"04",X"AF",X"21",X"D7",X"38",X"32",X"E7",X"49",X"11",
		X"E9",X"49",X"06",X"02",X"CD",X"54",X"3D",X"21",X"30",X"48",X"CD",X"00",X"03",X"79",X"32",X"E0",
		X"49",X"C3",X"EA",X"36",X"00",X"01",X"00",X"05",X"04",X"10",X"10",X"05",X"40",X"1D",X"FF",X"14",
		X"15",X"12",X"11",X"16",X"13",X"FF",X"AF",X"18",X"02",X"3E",X"01",X"32",X"01",X"50",X"32",X"05",
		X"50",X"32",X"06",X"50",X"C9",X"21",X"D1",X"40",X"01",X"14",X"03",X"3E",X"00",X"1E",X"00",X"CD",
		X"31",X"3D",X"DD",X"21",X"7E",X"3B",X"3A",X"01",X"48",X"CB",X"6F",X"28",X"04",X"DD",X"21",X"97",
		X"3B",X"CD",X"B2",X"3C",X"C9",X"DD",X"21",X"BB",X"3B",X"CD",X"B2",X"3C",X"DD",X"21",X"C7",X"3B",
		X"3A",X"01",X"48",X"CB",X"6F",X"28",X"04",X"DD",X"21",X"D6",X"3B",X"CD",X"B2",X"3C",X"3A",X"1B",
		X"48",X"E6",X"0C",X"C8",X"3A",X"E5",X"49",X"FE",X"02",X"C8",X"DD",X"21",X"E5",X"3B",X"CD",X"B2",
		X"3C",X"CD",X"A6",X"3E",X"E5",X"DD",X"E1",X"21",X"AC",X"41",X"1E",X"0D",X"06",X"06",X"0E",X"00",
		X"CD",X"8A",X"3D",X"C9",X"3A",X"1B",X"48",X"E6",X"03",X"21",X"71",X"39",X"07",X"06",X"00",X"4F",
		X"09",X"3A",X"01",X"48",X"CB",X"6F",X"28",X"01",X"23",X"7E",X"32",X"03",X"50",X"32",X"21",X"48",
		X"C9",X"00",X"01",X"00",X"00",X"01",X"00",X"01",X"01",X"3A",X"1B",X"48",X"E6",X"C0",X"07",X"07",
		X"21",X"8C",X"39",X"06",X"00",X"4F",X"09",X"7E",X"32",X"05",X"48",X"C9",X"00",X"01",X"02",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",
		X"5A",X"00",X"03",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"88",X"4B",X"06",X"28",X"CF",X"21",X"00",X"40",X"01",X"20",X"20",X"3E",X"00",X"1E",X"00",
		X"CD",X"99",X"3C",X"21",X"40",X"40",X"01",X"1C",X"01",X"3E",X"00",X"1E",X"0A",X"CD",X"31",X"3D",
		X"21",X"5F",X"40",X"01",X"1C",X"01",X"3E",X"00",X"1E",X"0A",X"CD",X"31",X"3D",X"C9",X"21",X"88",
		X"4B",X"06",X"28",X"CF",X"21",X"41",X"40",X"01",X"1C",X"1E",X"3E",X"00",X"1E",X"00",X"CD",X"99",
		X"3C",X"C9",X"21",X"BF",X"40",X"DD",X"21",X"0F",X"48",X"1E",X"0A",X"06",X"06",X"0E",X"00",X"CD",
		X"8A",X"3D",X"21",X"FF",X"42",X"DD",X"21",X"15",X"48",X"1E",X"0A",X"06",X"06",X"0E",X"00",X"CD",
		X"8A",X"3D",X"21",X"DF",X"41",X"DD",X"21",X"09",X"48",X"1E",X"0A",X"06",X"06",X"0E",X"00",X"CD",
		X"8A",X"3D",X"C9",X"DD",X"21",X"45",X"3A",X"06",X"0B",X"C5",X"DD",X"6E",X"00",X"DD",X"66",X"01",
		X"DD",X"7E",X"02",X"DD",X"5E",X"03",X"01",X"02",X"02",X"CD",X"1E",X"3D",X"01",X"04",X"00",X"DD",
		X"09",X"C1",X"10",X"E5",X"C9",X"B9",X"40",X"E0",X"11",X"F9",X"40",X"E4",X"12",X"39",X"41",X"E8",
		X"13",X"79",X"41",X"DC",X"11",X"B9",X"41",X"E0",X"13",X"F9",X"41",X"E4",X"12",X"39",X"42",X"E8",
		X"15",X"79",X"42",X"00",X"00",X"B9",X"42",X"EC",X"11",X"F9",X"42",X"E4",X"16",X"39",X"43",X"F0",
		X"12",X"DD",X"21",X"79",X"3A",X"CD",X"B2",X"3C",X"C9",X"00",X"02",X"7F",X"40",X"00",X"0D",X"31",
		X"50",X"02",X"9F",X"41",X"00",X"0D",X"48",X"49",X"02",X"BF",X"42",X"00",X"0D",X"32",X"50",X"00",
		X"00",X"14",X"CF",X"40",X"00",X"0B",X"50",X"55",X"53",X"48",X"20",X"31",X"20",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",X"00",X"15",X"CD",X"40",X"00",
		X"0C",X"50",X"55",X"53",X"48",X"20",X"32",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"20",
		X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",X"00",X"09",X"6F",X"41",X"00",X"0B",X"4D",X"4F",X"52",
		X"45",X"20",X"43",X"4F",X"49",X"4E",X"00",X"00",X"13",X"CD",X"40",X"00",X"0E",X"32",X"20",X"50",
		X"4C",X"41",X"59",X"45",X"52",X"53",X"20",X"4D",X"4F",X"52",X"45",X"20",X"43",X"4F",X"49",X"4E",
		X"00",X"00",X"0F",X"22",X"41",X"00",X"0A",X"40",X"20",X"31",X"39",X"38",X"33",X"20",X"53",X"41",
		X"4E",X"52",X"49",X"54",X"53",X"55",X"00",X"00",X"06",X"69",X"41",X"00",X"0A",X"43",X"52",X"45",
		X"44",X"49",X"54",X"00",X"00",X"02",X"E0",X"40",X"00",X"0C",X"4C",X"3D",X"00",X"25",X"3B",X"3B",
		X"3B",X"51",X"3B",X"67",X"3B",X"00",X"0F",X"26",X"41",X"00",X"0D",X"31",X"20",X"43",X"4F",X"49",
		X"4E",X"20",X"31",X"20",X"43",X"52",X"45",X"44",X"49",X"54",X"00",X"00",X"0F",X"26",X"41",X"00",
		X"0D",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"32",X"20",X"43",X"52",X"45",X"44",X"49",X"54",
		X"00",X"00",X"0F",X"26",X"41",X"00",X"0D",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"33",X"20",
		X"43",X"52",X"45",X"44",X"49",X"54",X"00",X"00",X"10",X"26",X"41",X"00",X"0D",X"32",X"20",X"43",
		X"4F",X"49",X"4E",X"53",X"20",X"31",X"20",X"43",X"52",X"45",X"44",X"49",X"54",X"00",X"00",X"12",
		X"F2",X"40",X"00",X"06",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"20",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"5F",X"31",X"00",X"00",X"12",X"F2",X"40",X"00",X"06",X"47",X"41",X"4D",
		X"45",X"20",X"4F",X"56",X"45",X"52",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"5F",X"32",X"00",
		X"00",X"04",X"A0",X"41",X"00",X"0A",X"54",X"49",X"4D",X"45",X"00",X"00",X"05",X"B2",X"41",X"00",
		X"0A",X"52",X"45",X"41",X"44",X"59",X"00",X"00",X"08",X"8F",X"41",X"00",X"0A",X"50",X"4C",X"41",
		X"59",X"45",X"52",X"20",X"31",X"00",X"00",X"08",X"8F",X"41",X"00",X"0A",X"50",X"4C",X"41",X"59",
		X"45",X"52",X"20",X"32",X"00",X"00",X"13",X"EC",X"40",X"00",X"0A",X"45",X"58",X"54",X"52",X"41",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"08",X"0F",X"00",X"07",X"08",X"04",X"00",X"07",X"08",X"01",X"00",
		X"07",X"08",X"03",X"00",X"03",X"08",X"05",X"00",X"03",X"02",X"07",X"00",X"07",X"08",X"05",X"00",
		X"07",X"0C",X"00",X"00",X"07",X"03",X"05",X"0D",X"00",X"00",X"07",X"0D",X"07",X"01",X"05",X"0D",
		X"03",X"05",X"02",X"0D",X"08",X"09",X"06",X"0D",X"02",X"05",X"08",X"0D",X"01",X"04",X"03",X"00",
		X"04",X"0A",X"05",X"00",X"01",X"03",X"00",X"00",X"05",X"08",X"00",X"00",X"03",X"02",X"00",X"00",
		X"07",X"08",X"01",X"00",X"03",X"01",X"07",X"00",X"02",X"03",X"00",X"00",X"09",X"0E",X"02",X"00",
		X"05",X"03",X"08",X"00",X"00",X"00",X"00",X"00",X"03",X"05",X"0F",X"00",X"03",X"0D",X"07",X"00",
		X"01",X"0D",X"07",X"00",X"0F",X"0D",X"07",X"0D",X"01",X"03",X"0E",X"00",X"05",X"0D",X"07",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5F",X"73",X"23",X"0B",X"79",X"B0",X"20",X"F9",X"C9",X"C5",X"E5",X"77",X"CD",X"43",X"3D",X"23",
		X"10",X"F9",X"F5",X"3E",X"23",X"06",X"01",X"FF",X"F1",X"E1",X"CD",X"4D",X"3D",X"C1",X"0D",X"20",
		X"E8",X"C9",X"DD",X"4E",X"00",X"DD",X"23",X"DD",X"7E",X"00",X"B7",X"C8",X"47",X"DD",X"23",X"DD",
		X"6E",X"00",X"DD",X"23",X"DD",X"66",X"00",X"DD",X"23",X"DD",X"7E",X"00",X"DD",X"23",X"B7",X"20",
		X"11",X"DD",X"5E",X"00",X"DD",X"23",X"DD",X"7E",X"00",X"CD",X"F3",X"3C",X"DD",X"23",X"10",X"F6",
		X"18",X"D5",X"DD",X"7E",X"00",X"DD",X"5E",X"01",X"CD",X"F3",X"3C",X"DD",X"23",X"DD",X"23",X"10",
		X"F1",X"18",X"C4",X"77",X"CD",X"43",X"3D",X"CD",X"4D",X"3D",X"79",X"B7",X"C8",X"C5",X"3E",X"23",
		X"41",X"FF",X"C1",X"C9",X"C5",X"E5",X"DD",X"7E",X"00",X"B7",X"28",X"04",X"77",X"CD",X"43",X"3D",
		X"DD",X"23",X"23",X"10",X"F1",X"E1",X"CD",X"4D",X"3D",X"C1",X"0D",X"20",X"E7",X"C9",X"C5",X"E5",
		X"77",X"CD",X"43",X"3D",X"23",X"3C",X"10",X"F8",X"E1",X"CD",X"4D",X"3D",X"C1",X"0D",X"20",X"EE",
		X"C9",X"C5",X"E5",X"77",X"CD",X"43",X"3D",X"23",X"10",X"F9",X"E1",X"CD",X"4D",X"3D",X"C1",X"0D",
		X"20",X"EF",X"C9",X"E5",X"D5",X"11",X"00",X"04",X"19",X"D1",X"73",X"E1",X"C9",X"D5",X"11",X"20",
		X"00",X"19",X"D1",X"C9",X"B7",X"1A",X"8E",X"FE",X"0A",X"38",X"02",X"D6",X"0A",X"12",X"3F",X"1B",
		X"2B",X"10",X"F2",X"C9",X"B7",X"1A",X"9E",X"30",X"02",X"C6",X"0A",X"12",X"1B",X"2B",X"10",X"F5",
		X"C9",X"1A",X"BE",X"38",X"08",X"20",X"09",X"13",X"23",X"10",X"F6",X"AF",X"C9",X"3E",X"01",X"C9",
		X"3E",X"02",X"C9",X"78",X"85",X"6F",X"79",X"84",X"67",X"C9",X"DD",X"7E",X"00",X"05",X"28",X"08",
		X"FE",X"00",X"20",X"03",X"B9",X"28",X"03",X"0D",X"C6",X"30",X"77",X"CD",X"43",X"3D",X"CD",X"4D",
		X"3D",X"DD",X"23",X"78",X"B7",X"20",X"E3",X"C9",X"7E",X"FE",X"FF",X"C8",X"FF",X"23",X"18",X"F8",
		X"7E",X"FE",X"FF",X"C8",X"23",X"4E",X"23",X"46",X"23",X"FF",X"18",X"F4",X"7D",X"FE",X"00",X"20",
		X"02",X"3E",X"FF",X"ED",X"44",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"5F",X"7C",X"ED",X"44",X"C6",
		X"10",X"ED",X"44",X"E6",X"F8",X"6F",X"26",X"00",X"54",X"29",X"29",X"19",X"11",X"00",X"40",X"19",
		X"C9",X"CB",X"27",X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"C9",X"0E",X"01",X"B7",X"28",X"05",
		X"3D",X"CB",X"21",X"18",X"F8",X"79",X"C9",X"06",X"04",X"0E",X"00",X"CB",X"3F",X"38",X"03",X"0C",
		X"10",X"F9",X"79",X"C9",X"3A",X"01",X"48",X"CB",X"7F",X"C8",X"DD",X"21",X"0F",X"48",X"11",X"14",
		X"48",X"01",X"BF",X"40",X"CB",X"6F",X"3E",X"0A",X"28",X"0C",X"DD",X"21",X"15",X"48",X"11",X"1A",
		X"48",X"01",X"FF",X"42",X"3E",X"0A",X"F5",X"C5",X"06",X"06",X"CD",X"54",X"3D",X"E1",X"F1",X"06",
		X"06",X"5F",X"0E",X"00",X"CD",X"8A",X"3D",X"3A",X"01",X"48",X"11",X"0F",X"48",X"CB",X"6F",X"28",
		X"03",X"11",X"15",X"48",X"06",X"06",X"D5",X"21",X"09",X"48",X"CD",X"71",X"3D",X"E1",X"FE",X"02",
		X"20",X"18",X"11",X"09",X"48",X"01",X"06",X"00",X"ED",X"B0",X"DD",X"21",X"09",X"48",X"21",X"DF",
		X"41",X"06",X"06",X"1E",X"0A",X"0E",X"00",X"CD",X"8A",X"3D",X"3A",X"1B",X"48",X"E6",X"0C",X"FE",
		X"00",X"C8",X"3A",X"E5",X"49",X"FE",X"02",X"C8",X"CD",X"A6",X"3E",X"3A",X"01",X"48",X"11",X"0F",
		X"48",X"CB",X"6F",X"28",X"03",X"11",X"15",X"48",X"06",X"06",X"CD",X"71",X"3D",X"FE",X"01",X"C8",
		X"3E",X"0E",X"16",X"00",X"5A",X"CD",X"20",X"2C",X"21",X"E5",X"49",X"34",X"21",X"E6",X"49",X"34",
		X"46",X"05",X"CD",X"EF",X"3E",X"C9",X"21",X"C5",X"3E",X"3A",X"1B",X"48",X"E6",X"0C",X"CB",X"3F",
		X"CB",X"3F",X"3D",X"CD",X"E1",X"3D",X"EB",X"3A",X"E5",X"49",X"CB",X"27",X"5F",X"CB",X"27",X"83",
		X"5F",X"16",X"00",X"19",X"C9",X"CB",X"3E",X"D7",X"3E",X"E3",X"3E",X"00",X"02",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"01",X"04",X"00",
		X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"C5",
		X"21",X"40",X"40",X"1E",X"1E",X"01",X"01",X"01",X"3E",X"2D",X"CD",X"31",X"3D",X"1E",X"0A",X"3E",
		X"3D",X"01",X"01",X"01",X"CD",X"31",X"3D",X"C1",X"78",X"F6",X"30",X"01",X"01",X"01",X"CD",X"31",
		X"3D",X"C9",X"21",X"60",X"43",X"3A",X"E1",X"49",X"FE",X"08",X"38",X"0B",X"D6",X"08",X"F5",X"3E",
		X"FF",X"CD",X"29",X"3F",X"F1",X"18",X"F1",X"C6",X"F7",X"47",X"1E",X"0B",X"3A",X"DA",X"49",X"CB",
		X"47",X"28",X"02",X"1E",X"0F",X"78",X"01",X"01",X"01",X"CD",X"31",X"3D",X"11",X"C0",X"FF",X"19",
		X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"31",X"B0",X"4D",X"21",X"50",X"4B",X"06",X"20",
		X"CF",X"3E",X"23",X"06",X"01",X"FF",X"FD",X"21",X"50",X"4B",X"06",X"08",X"C5",X"FD",X"7E",X"00",
		X"FD",X"B6",X"01",X"28",X"03",X"CD",X"73",X"3F",X"01",X"04",X"00",X"FD",X"09",X"C1",X"10",X"EC",
		X"C3",X"51",X"3F",X"FD",X"7E",X"02",X"B7",X"28",X"04",X"FD",X"35",X"02",X"C9",X"FD",X"36",X"02",
		X"08",X"FD",X"7E",X"03",X"3C",X"FD",X"77",X"03",X"FE",X"20",X"28",X"14",X"FD",X"66",X"00",X"FD",
		X"6E",X"01",X"CD",X"BC",X"3D",X"3E",X"10",X"1E",X"10",X"01",X"02",X"02",X"CD",X"1E",X"3D",X"C9",
		X"FD",X"66",X"00",X"FD",X"6E",X"01",X"E5",X"CD",X"9E",X"0F",X"7E",X"E6",X"0F",X"77",X"E1",X"F5",
		X"CD",X"BC",X"3D",X"F1",X"1E",X"01",X"DD",X"21",X"77",X"89",X"CD",X"50",X"89",X"FD",X"E5",X"E1",
		X"06",X"04",X"CF",X"C9",X"FD",X"E5",X"FD",X"21",X"50",X"4B",X"06",X"08",X"FD",X"7E",X"00",X"FD",
		X"B6",X"01",X"28",X"16",X"FD",X"7E",X"00",X"BC",X"20",X"06",X"FD",X"7E",X"01",X"BD",X"28",X"07",
		X"11",X"04",X"00",X"FD",X"19",X"10",X"E5",X"37",X"18",X"11",X"E5",X"CD",X"9E",X"0F",X"E6",X"0F",
		X"F6",X"80",X"77",X"E1",X"FD",X"74",X"00",X"FD",X"75",X"01",X"A7",X"FD",X"E1",X"C9",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
